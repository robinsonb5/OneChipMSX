-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b0bb4",
     9 => x"bc080b0b",
    10 => x"0bb4c008",
    11 => x"0b0b0bb4",
    12 => x"c4080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"b4c40c0b",
    16 => x"0b0bb4c0",
    17 => x"0c0b0b0b",
    18 => x"b4bc0c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0baad4",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"b4bc70b9",
    57 => x"f4278b38",
    58 => x"80717084",
    59 => x"05530c81",
    60 => x"e2048c51",
    61 => x"8bb00402",
    62 => x"fc050df8",
    63 => x"80518f0b",
    64 => x"b4cc0c9f",
    65 => x"0bb4d00c",
    66 => x"a0717081",
    67 => x"055334b4",
    68 => x"d008ff05",
    69 => x"b4d00cb4",
    70 => x"d0088025",
    71 => x"eb38b4cc",
    72 => x"08ff05b4",
    73 => x"cc0cb4cc",
    74 => x"088025d7",
    75 => x"38028405",
    76 => x"0d0402f0",
    77 => x"050df880",
    78 => x"53f8a054",
    79 => x"83bf5273",
    80 => x"70810555",
    81 => x"33517073",
    82 => x"70810555",
    83 => x"34ff1252",
    84 => x"718025eb",
    85 => x"38fbc053",
    86 => x"9f52a073",
    87 => x"70810555",
    88 => x"34ff1252",
    89 => x"718025f2",
    90 => x"38029005",
    91 => x"0d0402f4",
    92 => x"050d7453",
    93 => x"8e0bb4cc",
    94 => x"08258f38",
    95 => x"82b22db4",
    96 => x"cc08ff05",
    97 => x"b4cc0c82",
    98 => x"f404b4cc",
    99 => x"08b4d008",
   100 => x"5351728a",
   101 => x"2e098106",
   102 => x"b7387151",
   103 => x"719f24a0",
   104 => x"38b4cc08",
   105 => x"a02911f8",
   106 => x"80115151",
   107 => x"a07134b4",
   108 => x"d0088105",
   109 => x"b4d00cb4",
   110 => x"d008519f",
   111 => x"7125e238",
   112 => x"800bb4d0",
   113 => x"0cb4cc08",
   114 => x"8105b4cc",
   115 => x"0c83e404",
   116 => x"70a02912",
   117 => x"f8801151",
   118 => x"51727134",
   119 => x"b4d00881",
   120 => x"05b4d00c",
   121 => x"b4d008a0",
   122 => x"2e098106",
   123 => x"8e38800b",
   124 => x"b4d00cb4",
   125 => x"cc088105",
   126 => x"b4cc0c02",
   127 => x"8c050d04",
   128 => x"02e8050d",
   129 => x"77795656",
   130 => x"880bfc16",
   131 => x"77712c8f",
   132 => x"06545254",
   133 => x"80537272",
   134 => x"25953871",
   135 => x"53fbe014",
   136 => x"51877134",
   137 => x"8114ff14",
   138 => x"545472f1",
   139 => x"387153f9",
   140 => x"1576712c",
   141 => x"87065351",
   142 => x"71802e8b",
   143 => x"38fbe014",
   144 => x"51717134",
   145 => x"81145472",
   146 => x"8e249538",
   147 => x"8f733153",
   148 => x"fbe01451",
   149 => x"a0713481",
   150 => x"14ff1454",
   151 => x"5472f138",
   152 => x"0298050d",
   153 => x"0402ec05",
   154 => x"0d800bb4",
   155 => x"d40cf68c",
   156 => x"08f69008",
   157 => x"71882c56",
   158 => x"5481ff06",
   159 => x"52737225",
   160 => x"88387154",
   161 => x"820bb4d4",
   162 => x"0c72882c",
   163 => x"7381ff06",
   164 => x"54557473",
   165 => x"258b3872",
   166 => x"b4d40884",
   167 => x"07b4d40c",
   168 => x"5573842b",
   169 => x"86a07125",
   170 => x"83713170",
   171 => x"0b0b0bb1",
   172 => x"a40c8171",
   173 => x"2bff05f6",
   174 => x"880cfecc",
   175 => x"13ff122c",
   176 => x"788829ff",
   177 => x"94057081",
   178 => x"2cb4d408",
   179 => x"52585255",
   180 => x"51525476",
   181 => x"802e8538",
   182 => x"70810751",
   183 => x"70f6940c",
   184 => x"71098105",
   185 => x"f6800c72",
   186 => x"098105f6",
   187 => x"840c0294",
   188 => x"050d0402",
   189 => x"f4050d74",
   190 => x"53727081",
   191 => x"055480f5",
   192 => x"2d527180",
   193 => x"2e893871",
   194 => x"5182ee2d",
   195 => x"85f90402",
   196 => x"8c050d04",
   197 => x"02f8050d",
   198 => x"a28d2d80",
   199 => x"da51a3c4",
   200 => x"2db4bc08",
   201 => x"812a7081",
   202 => x"06515271",
   203 => x"802ee938",
   204 => x"0288050d",
   205 => x"0402f405",
   206 => x"0db9e408",
   207 => x"99c406b3",
   208 => x"940b80f5",
   209 => x"2d525270",
   210 => x"802e8638",
   211 => x"71848007",
   212 => x"52b2cc0b",
   213 => x"80f52d72",
   214 => x"07b2e40b",
   215 => x"80f52d70",
   216 => x"812a7081",
   217 => x"06515354",
   218 => x"5270802e",
   219 => x"86387182",
   220 => x"80075272",
   221 => x"81065170",
   222 => x"802e8538",
   223 => x"71880752",
   224 => x"b2f00b80",
   225 => x"f52d7084",
   226 => x"2b730781",
   227 => x"8432b4bc",
   228 => x"0c51028c",
   229 => x"050d0402",
   230 => x"f4050d74",
   231 => x"70818432",
   232 => x"b9e40c70",
   233 => x"83065253",
   234 => x"70b2c40b",
   235 => x"880581b7",
   236 => x"2d72892a",
   237 => x"70810651",
   238 => x"5170b394",
   239 => x"0b81b72d",
   240 => x"72832a81",
   241 => x"0673882a",
   242 => x"70810651",
   243 => x"52527080",
   244 => x"2e853871",
   245 => x"82075271",
   246 => x"b2e40b81",
   247 => x"b72d7284",
   248 => x"2c708306",
   249 => x"515170b2",
   250 => x"f00b81b7",
   251 => x"2d70b4bc",
   252 => x"0c028c05",
   253 => x"0d0402d4",
   254 => x"050dadd8",
   255 => x"5185f32d",
   256 => x"9bb92db4",
   257 => x"bc08802e",
   258 => x"82ab3886",
   259 => x"b52db4bc",
   260 => x"08538ea8",
   261 => x"2db4bc08",
   262 => x"54b4bc08",
   263 => x"802e8297",
   264 => x"389df42d",
   265 => x"b4bc0880",
   266 => x"2e8738ad",
   267 => x"f05188be",
   268 => x"0497a52d",
   269 => x"b4bc0880",
   270 => x"2e9c38ae",
   271 => x"b05185f3",
   272 => x"2d86942d",
   273 => x"72840753",
   274 => x"810bfec4",
   275 => x"0c72fec0",
   276 => x"0c725187",
   277 => x"972d840b",
   278 => x"fec40cae",
   279 => x"f85185f3",
   280 => x"2daf9052",
   281 => x"b4dc5194",
   282 => x"ba2db4bc",
   283 => x"089838af",
   284 => x"9c5185f3",
   285 => x"2dafb452",
   286 => x"b4dc5194",
   287 => x"ba2db4bc",
   288 => x"08802e81",
   289 => x"b038afc0",
   290 => x"5185f32d",
   291 => x"b4e00857",
   292 => x"8077595a",
   293 => x"767a2e8b",
   294 => x"38811a78",
   295 => x"812a595a",
   296 => x"77f738f7",
   297 => x"1a5a8077",
   298 => x"25818038",
   299 => x"79527751",
   300 => x"84802db4",
   301 => x"e852b4dc",
   302 => x"5196ff2d",
   303 => x"b4bc0853",
   304 => x"b4bc0880",
   305 => x"2e80c938",
   306 => x"b4e85b80",
   307 => x"5989fd04",
   308 => x"7a708405",
   309 => x"5c087081",
   310 => x"ff067188",
   311 => x"2c7081ff",
   312 => x"0673902c",
   313 => x"7081ff06",
   314 => x"75982afe",
   315 => x"c80cfec8",
   316 => x"0c58fec8",
   317 => x"0c57fec8",
   318 => x"0c841a5a",
   319 => x"53765384",
   320 => x"80772584",
   321 => x"38848053",
   322 => x"727924c4",
   323 => x"388a9b04",
   324 => x"afdc5185",
   325 => x"f32d7254",
   326 => x"8ab704b4",
   327 => x"dc5196d2",
   328 => x"2dfc8017",
   329 => x"81195957",
   330 => x"89a60482",
   331 => x"0bfec40c",
   332 => x"81548ab7",
   333 => x"04805473",
   334 => x"b4bc0c02",
   335 => x"ac050d04",
   336 => x"02f8050d",
   337 => x"a4942d81",
   338 => x"f72d8151",
   339 => x"84e52dfe",
   340 => x"c4528172",
   341 => x"0ca1d42d",
   342 => x"a1d42d84",
   343 => x"720c87f6",
   344 => x"2db1a851",
   345 => x"a5f22d80",
   346 => x"5184e52d",
   347 => x"0288050d",
   348 => x"0402f405",
   349 => x"0db1fc0b",
   350 => x"881180f5",
   351 => x"2d8c1288",
   352 => x"1180f52d",
   353 => x"70842b73",
   354 => x"078c1388",
   355 => x"1180f52d",
   356 => x"70882b73",
   357 => x"07941380",
   358 => x"f52d708c",
   359 => x"2b7207b4",
   360 => x"bc0c5353",
   361 => x"53535356",
   362 => x"52535102",
   363 => x"8c050d04",
   364 => x"02ec050d",
   365 => x"8cb85187",
   366 => x"972d810b",
   367 => x"fec40c8c",
   368 => x"b80bfec0",
   369 => x"0c840bfe",
   370 => x"c40c830b",
   371 => x"fecc0ca1",
   372 => x"ef2da488",
   373 => x"2da1d42d",
   374 => x"a1d42d81",
   375 => x"f72d8151",
   376 => x"84e52da1",
   377 => x"d42da1d4",
   378 => x"2d815184",
   379 => x"e52d87f6",
   380 => x"2db4bc08",
   381 => x"802e81dd",
   382 => x"38805184",
   383 => x"e52db1a8",
   384 => x"51a5f22d",
   385 => x"b9cc0809",
   386 => x"708306fe",
   387 => x"cc0c52b9",
   388 => x"c4088938",
   389 => x"b9c80880",
   390 => x"2e80e238",
   391 => x"fed00870",
   392 => x"81065152",
   393 => x"71802e80",
   394 => x"d438a48e",
   395 => x"2db9c408",
   396 => x"70b9c808",
   397 => x"70575556",
   398 => x"5280ff72",
   399 => x"25843880",
   400 => x"ff5280ff",
   401 => x"73258438",
   402 => x"80ff5371",
   403 => x"ff802584",
   404 => x"38ff8052",
   405 => x"72ff8025",
   406 => x"8438ff80",
   407 => x"53747231",
   408 => x"b9c40c73",
   409 => x"7331b9c8",
   410 => x"0ca4882d",
   411 => x"71882b83",
   412 => x"fe800673",
   413 => x"81ff0671",
   414 => x"07fed00c",
   415 => x"52a28d2d",
   416 => x"a6822db4",
   417 => x"bc085386",
   418 => x"b52db4bc",
   419 => x"08fec00c",
   420 => x"8af12db4",
   421 => x"bc08fed4",
   422 => x"0c86b52d",
   423 => x"b4bc08b4",
   424 => x"d8082e9c",
   425 => x"38b4bc08",
   426 => x"b4d80c84",
   427 => x"52725184",
   428 => x"e52da1d4",
   429 => x"2da1d42d",
   430 => x"ff125271",
   431 => x"8025ee38",
   432 => x"72802e89",
   433 => x"388a0bfe",
   434 => x"c40c8c84",
   435 => x"04820bfe",
   436 => x"c40c8c84",
   437 => x"04aff051",
   438 => x"85f32d82",
   439 => x"0bfec40c",
   440 => x"800bb4bc",
   441 => x"0c029405",
   442 => x"0d0402e8",
   443 => x"050d7779",
   444 => x"7b585555",
   445 => x"80537276",
   446 => x"25a33874",
   447 => x"70810556",
   448 => x"80f52d74",
   449 => x"70810556",
   450 => x"80f52d52",
   451 => x"5271712e",
   452 => x"86388151",
   453 => x"8e9f0481",
   454 => x"13538df6",
   455 => x"04805170",
   456 => x"b4bc0c02",
   457 => x"98050d04",
   458 => x"02d8050d",
   459 => x"800bb8f0",
   460 => x"0cb4e852",
   461 => x"80519cd9",
   462 => x"2db4bc08",
   463 => x"54b4bc08",
   464 => x"8c38b088",
   465 => x"5185f32d",
   466 => x"735593c3",
   467 => x"04805681",
   468 => x"0bb9940c",
   469 => x"8853b09c",
   470 => x"52b59e51",
   471 => x"8dea2db4",
   472 => x"bc08762e",
   473 => x"09810687",
   474 => x"38b4bc08",
   475 => x"b9940c88",
   476 => x"53b0a852",
   477 => x"b5ba518d",
   478 => x"ea2db4bc",
   479 => x"088738b4",
   480 => x"bc08b994",
   481 => x"0cb99408",
   482 => x"802e80f6",
   483 => x"38b8ae0b",
   484 => x"80f52db8",
   485 => x"af0b80f5",
   486 => x"2d71982b",
   487 => x"71902b07",
   488 => x"b8b00b80",
   489 => x"f52d7088",
   490 => x"2b7207b8",
   491 => x"b10b80f5",
   492 => x"2d7107b8",
   493 => x"e60b80f5",
   494 => x"2db8e70b",
   495 => x"80f52d71",
   496 => x"882b0753",
   497 => x"5f54525a",
   498 => x"56575573",
   499 => x"81abaa2e",
   500 => x"0981068d",
   501 => x"3875519d",
   502 => x"fb2db4bc",
   503 => x"08568fee",
   504 => x"047382d4",
   505 => x"d52e8738",
   506 => x"b0b45190",
   507 => x"af04b4e8",
   508 => x"5275519c",
   509 => x"d92db4bc",
   510 => x"0855b4bc",
   511 => x"08802e83",
   512 => x"c2388853",
   513 => x"b0a852b5",
   514 => x"ba518dea",
   515 => x"2db4bc08",
   516 => x"8938810b",
   517 => x"b8f00c90",
   518 => x"b5048853",
   519 => x"b09c52b5",
   520 => x"9e518dea",
   521 => x"2db4bc08",
   522 => x"802e8a38",
   523 => x"b0c85185",
   524 => x"f32d918f",
   525 => x"04b8e60b",
   526 => x"80f52d54",
   527 => x"7380d52e",
   528 => x"09810680",
   529 => x"ca38b8e7",
   530 => x"0b80f52d",
   531 => x"547381aa",
   532 => x"2e098106",
   533 => x"ba38800b",
   534 => x"b4e80b80",
   535 => x"f52d5654",
   536 => x"7481e92e",
   537 => x"83388154",
   538 => x"7481eb2e",
   539 => x"8c388055",
   540 => x"73752e09",
   541 => x"810682cb",
   542 => x"38b4f30b",
   543 => x"80f52d55",
   544 => x"748d38b4",
   545 => x"f40b80f5",
   546 => x"2d547382",
   547 => x"2e863880",
   548 => x"5593c304",
   549 => x"b4f50b80",
   550 => x"f52d70b8",
   551 => x"e80cff05",
   552 => x"b8ec0cb4",
   553 => x"f60b80f5",
   554 => x"2db4f70b",
   555 => x"80f52d58",
   556 => x"76057782",
   557 => x"80290570",
   558 => x"b8f40cb4",
   559 => x"f80b80f5",
   560 => x"2d70b988",
   561 => x"0cb8f008",
   562 => x"59575876",
   563 => x"802e81a3",
   564 => x"388853b0",
   565 => x"a852b5ba",
   566 => x"518dea2d",
   567 => x"b4bc0881",
   568 => x"e238b8e8",
   569 => x"0870842b",
   570 => x"b98c0c70",
   571 => x"b9840cb5",
   572 => x"8d0b80f5",
   573 => x"2db58c0b",
   574 => x"80f52d71",
   575 => x"82802905",
   576 => x"b58e0b80",
   577 => x"f52d7084",
   578 => x"80802912",
   579 => x"b58f0b80",
   580 => x"f52d7081",
   581 => x"800a2912",
   582 => x"70b9900c",
   583 => x"b9880871",
   584 => x"29b8f408",
   585 => x"0570b8f8",
   586 => x"0cb5950b",
   587 => x"80f52db5",
   588 => x"940b80f5",
   589 => x"2d718280",
   590 => x"2905b596",
   591 => x"0b80f52d",
   592 => x"70848080",
   593 => x"2912b597",
   594 => x"0b80f52d",
   595 => x"70982b81",
   596 => x"f00a0672",
   597 => x"0570b8fc",
   598 => x"0cfe117e",
   599 => x"297705b9",
   600 => x"800c5259",
   601 => x"5243545e",
   602 => x"51525952",
   603 => x"5d575957",
   604 => x"93c104b4",
   605 => x"fa0b80f5",
   606 => x"2db4f90b",
   607 => x"80f52d71",
   608 => x"82802905",
   609 => x"70b98c0c",
   610 => x"70a02983",
   611 => x"ff057089",
   612 => x"2a70b984",
   613 => x"0cb4ff0b",
   614 => x"80f52db4",
   615 => x"fe0b80f5",
   616 => x"2d718280",
   617 => x"290570b9",
   618 => x"900c7b71",
   619 => x"291e70b9",
   620 => x"800c7db8",
   621 => x"fc0c7305",
   622 => x"b8f80c55",
   623 => x"5e515155",
   624 => x"55815574",
   625 => x"b4bc0c02",
   626 => x"a8050d04",
   627 => x"02ec050d",
   628 => x"7670872c",
   629 => x"7180ff06",
   630 => x"555654b8",
   631 => x"f0088a38",
   632 => x"73882c74",
   633 => x"81ff0654",
   634 => x"55b4e852",
   635 => x"b8f40815",
   636 => x"519cd92d",
   637 => x"b4bc0854",
   638 => x"b4bc0880",
   639 => x"2eb338b8",
   640 => x"f008802e",
   641 => x"98387284",
   642 => x"29b4e805",
   643 => x"70085253",
   644 => x"9dfb2db4",
   645 => x"bc08f00a",
   646 => x"065394af",
   647 => x"047210b4",
   648 => x"e8057080",
   649 => x"e02d5253",
   650 => x"9eab2db4",
   651 => x"bc085372",
   652 => x"5473b4bc",
   653 => x"0c029405",
   654 => x"0d0402c8",
   655 => x"050d7f61",
   656 => x"5f5b800b",
   657 => x"b8fc08b9",
   658 => x"8008595d",
   659 => x"56b8f008",
   660 => x"762e8a38",
   661 => x"b8e80884",
   662 => x"2b5894e3",
   663 => x"04b98408",
   664 => x"842b5880",
   665 => x"59787827",
   666 => x"81a93878",
   667 => x"8f06a017",
   668 => x"5754738f",
   669 => x"38b4e852",
   670 => x"76518117",
   671 => x"579cd92d",
   672 => x"b4e85680",
   673 => x"7680f52d",
   674 => x"56547474",
   675 => x"2e833881",
   676 => x"547481e5",
   677 => x"2e80f638",
   678 => x"81707506",
   679 => x"555d7380",
   680 => x"2e80ea38",
   681 => x"8b1680f5",
   682 => x"2d98065a",
   683 => x"7980de38",
   684 => x"8b537d52",
   685 => x"75518dea",
   686 => x"2db4bc08",
   687 => x"80cf389c",
   688 => x"1608519d",
   689 => x"fb2db4bc",
   690 => x"08841c0c",
   691 => x"9a1680e0",
   692 => x"2d519eab",
   693 => x"2db4bc08",
   694 => x"b4bc0888",
   695 => x"1d0cb4bc",
   696 => x"085555b8",
   697 => x"f008802e",
   698 => x"98389416",
   699 => x"80e02d51",
   700 => x"9eab2db4",
   701 => x"bc08902b",
   702 => x"83fff00a",
   703 => x"06701651",
   704 => x"5473881c",
   705 => x"0c797b0c",
   706 => x"7c5496c9",
   707 => x"04811959",
   708 => x"94e504b8",
   709 => x"f008802e",
   710 => x"ae387b51",
   711 => x"93cc2db4",
   712 => x"bc08b4bc",
   713 => x"0880ffff",
   714 => x"fff80655",
   715 => x"5c7380ff",
   716 => x"fffff82e",
   717 => x"9238b4bc",
   718 => x"08fe05b8",
   719 => x"e80829b8",
   720 => x"f8080557",
   721 => x"94e30480",
   722 => x"5473b4bc",
   723 => x"0c02b805",
   724 => x"0d0402f4",
   725 => x"050d7470",
   726 => x"08810571",
   727 => x"0c7008b8",
   728 => x"ec080653",
   729 => x"53718e38",
   730 => x"88130851",
   731 => x"93cc2db4",
   732 => x"bc088814",
   733 => x"0c810bb4",
   734 => x"bc0c028c",
   735 => x"050d0402",
   736 => x"f0050d75",
   737 => x"881108fe",
   738 => x"05b8e808",
   739 => x"29b8f808",
   740 => x"117208b8",
   741 => x"ec080605",
   742 => x"79555354",
   743 => x"549cd92d",
   744 => x"0290050d",
   745 => x"04b8f008",
   746 => x"b4bc0c04",
   747 => x"02f4050d",
   748 => x"d45281ff",
   749 => x"720c7108",
   750 => x"5381ff72",
   751 => x"0c72882b",
   752 => x"83fe8006",
   753 => x"72087081",
   754 => x"ff065152",
   755 => x"5381ff72",
   756 => x"0c727107",
   757 => x"882b7208",
   758 => x"7081ff06",
   759 => x"51525381",
   760 => x"ff720c72",
   761 => x"7107882b",
   762 => x"72087081",
   763 => x"ff067207",
   764 => x"b4bc0c52",
   765 => x"53028c05",
   766 => x"0d0402f4",
   767 => x"050d7476",
   768 => x"7181ff06",
   769 => x"d40c5353",
   770 => x"b9980885",
   771 => x"3871892b",
   772 => x"5271982a",
   773 => x"d40c7190",
   774 => x"2a7081ff",
   775 => x"06d40c51",
   776 => x"71882a70",
   777 => x"81ff06d4",
   778 => x"0c517181",
   779 => x"ff06d40c",
   780 => x"72902a70",
   781 => x"81ff06d4",
   782 => x"0c51d408",
   783 => x"7081ff06",
   784 => x"515182b8",
   785 => x"bf527081",
   786 => x"ff2e0981",
   787 => x"06943881",
   788 => x"ff0bd40c",
   789 => x"d4087081",
   790 => x"ff06ff14",
   791 => x"54515171",
   792 => x"e53870b4",
   793 => x"bc0c028c",
   794 => x"050d0402",
   795 => x"fc050d81",
   796 => x"c75181ff",
   797 => x"0bd40cff",
   798 => x"11517080",
   799 => x"25f43802",
   800 => x"84050d04",
   801 => x"02f0050d",
   802 => x"98eb2d8f",
   803 => x"cf538052",
   804 => x"87fc80f7",
   805 => x"5197fa2d",
   806 => x"b4bc0854",
   807 => x"b4bc0881",
   808 => x"2e098106",
   809 => x"a33881ff",
   810 => x"0bd40c82",
   811 => x"0a52849c",
   812 => x"80e95197",
   813 => x"fa2db4bc",
   814 => x"088b3881",
   815 => x"ff0bd40c",
   816 => x"735399ce",
   817 => x"0498eb2d",
   818 => x"ff135372",
   819 => x"c13872b4",
   820 => x"bc0c0290",
   821 => x"050d0402",
   822 => x"f4050d81",
   823 => x"ff0bd40c",
   824 => x"93538052",
   825 => x"87fc80c1",
   826 => x"5197fa2d",
   827 => x"b4bc088b",
   828 => x"3881ff0b",
   829 => x"d40c8153",
   830 => x"9a840498",
   831 => x"eb2dff13",
   832 => x"5372df38",
   833 => x"72b4bc0c",
   834 => x"028c050d",
   835 => x"0402f005",
   836 => x"0d98eb2d",
   837 => x"83aa5284",
   838 => x"9c80c851",
   839 => x"97fa2db4",
   840 => x"bc08812e",
   841 => x"09810692",
   842 => x"3897ac2d",
   843 => x"b4bc0883",
   844 => x"ffff0653",
   845 => x"7283aa2e",
   846 => x"973899d7",
   847 => x"2d9acb04",
   848 => x"81549bb0",
   849 => x"04b0d451",
   850 => x"85f32d80",
   851 => x"549bb004",
   852 => x"81ff0bd4",
   853 => x"0cb15399",
   854 => x"842db4bc",
   855 => x"08802e80",
   856 => x"c0388052",
   857 => x"87fc80fa",
   858 => x"5197fa2d",
   859 => x"b4bc08b1",
   860 => x"3881ff0b",
   861 => x"d40cd408",
   862 => x"5381ff0b",
   863 => x"d40c81ff",
   864 => x"0bd40c81",
   865 => x"ff0bd40c",
   866 => x"81ff0bd4",
   867 => x"0c72862a",
   868 => x"708106b4",
   869 => x"bc085651",
   870 => x"5372802e",
   871 => x"93389ac0",
   872 => x"0472822e",
   873 => x"ff9f38ff",
   874 => x"135372ff",
   875 => x"aa387254",
   876 => x"73b4bc0c",
   877 => x"0290050d",
   878 => x"0402f405",
   879 => x"0d810bb9",
   880 => x"980cd008",
   881 => x"708f2a70",
   882 => x"81065151",
   883 => x"5372f338",
   884 => x"72d00c98",
   885 => x"eb2db0e4",
   886 => x"5185f32d",
   887 => x"d008708f",
   888 => x"2a708106",
   889 => x"51515372",
   890 => x"f338810b",
   891 => x"d00c80e3",
   892 => x"53805284",
   893 => x"d480c051",
   894 => x"97fa2db4",
   895 => x"bc08812e",
   896 => x"9a387282",
   897 => x"2e098106",
   898 => x"8c38b0f0",
   899 => x"5185f32d",
   900 => x"80539cd0",
   901 => x"04ff1353",
   902 => x"72d7389a",
   903 => x"8d2db4bc",
   904 => x"08b9980c",
   905 => x"b4bc088b",
   906 => x"38815287",
   907 => x"fc80d051",
   908 => x"97fa2d81",
   909 => x"ff0bd40c",
   910 => x"d008708f",
   911 => x"2a708106",
   912 => x"51515372",
   913 => x"f33872d0",
   914 => x"0c81ff0b",
   915 => x"d40c8153",
   916 => x"72b4bc0c",
   917 => x"028c050d",
   918 => x"0402e805",
   919 => x"0d785580",
   920 => x"5681ff0b",
   921 => x"d40cd008",
   922 => x"708f2a70",
   923 => x"81065151",
   924 => x"5372f338",
   925 => x"82810bd0",
   926 => x"0c81ff0b",
   927 => x"d40c7752",
   928 => x"87fc80d1",
   929 => x"5197fa2d",
   930 => x"80dbc6df",
   931 => x"54b4bc08",
   932 => x"802e8a38",
   933 => x"b1885185",
   934 => x"f32d9deb",
   935 => x"0481ff0b",
   936 => x"d40cd408",
   937 => x"7081ff06",
   938 => x"51537281",
   939 => x"fe2e0981",
   940 => x"069d3880",
   941 => x"ff5397ac",
   942 => x"2db4bc08",
   943 => x"75708405",
   944 => x"570cff13",
   945 => x"53728025",
   946 => x"ed388156",
   947 => x"9dd504ff",
   948 => x"145473c9",
   949 => x"3881ff0b",
   950 => x"d40cd008",
   951 => x"708f2a70",
   952 => x"81065151",
   953 => x"5372f338",
   954 => x"72d00c75",
   955 => x"b4bc0c02",
   956 => x"98050d04",
   957 => x"b99808b4",
   958 => x"bc0c0402",
   959 => x"f4050d74",
   960 => x"70882a83",
   961 => x"fe800670",
   962 => x"72982a07",
   963 => x"72882b87",
   964 => x"fc808006",
   965 => x"73982b81",
   966 => x"f00a0671",
   967 => x"730707b4",
   968 => x"bc0c5651",
   969 => x"5351028c",
   970 => x"050d0402",
   971 => x"f8050d02",
   972 => x"8e0580f5",
   973 => x"2d74882b",
   974 => x"077083ff",
   975 => x"ff06b4bc",
   976 => x"0c510288",
   977 => x"050d0402",
   978 => x"fc050d72",
   979 => x"5180710c",
   980 => x"800b8412",
   981 => x"0c028405",
   982 => x"0d0402f0",
   983 => x"050d7570",
   984 => x"08841208",
   985 => x"535353ff",
   986 => x"5471712e",
   987 => x"a838a48e",
   988 => x"2d841308",
   989 => x"70842914",
   990 => x"88117008",
   991 => x"7081ff06",
   992 => x"84180881",
   993 => x"11870684",
   994 => x"1a0c5351",
   995 => x"55515151",
   996 => x"a4882d71",
   997 => x"5473b4bc",
   998 => x"0c029005",
   999 => x"0d0402f0",
  1000 => x"050da48e",
  1001 => x"2de008e4",
  1002 => x"08718b2a",
  1003 => x"70810651",
  1004 => x"53555270",
  1005 => x"802e9d38",
  1006 => x"b99c0870",
  1007 => x"8429b9a4",
  1008 => x"057381ff",
  1009 => x"06710c51",
  1010 => x"51b99c08",
  1011 => x"81118706",
  1012 => x"b99c0c51",
  1013 => x"738b2a70",
  1014 => x"81065151",
  1015 => x"70802e81",
  1016 => x"8938b3ec",
  1017 => x"088429b9",
  1018 => x"d4057481",
  1019 => x"ff06710c",
  1020 => x"51b3ec08",
  1021 => x"8105b3ec",
  1022 => x"0c850bb3",
  1023 => x"e80cb3ec",
  1024 => x"08b3e408",
  1025 => x"2e098106",
  1026 => x"81863880",
  1027 => x"0bb3ec0c",
  1028 => x"b9d40870",
  1029 => x"8306b9cc",
  1030 => x"0c70852a",
  1031 => x"708106b9",
  1032 => x"c8085651",
  1033 => x"52527080",
  1034 => x"2e8e38b9",
  1035 => x"dc08fe80",
  1036 => x"3213b9c8",
  1037 => x"0ca0bf04",
  1038 => x"b9dc0813",
  1039 => x"b9c80c71",
  1040 => x"842a7081",
  1041 => x"06b9c408",
  1042 => x"54515170",
  1043 => x"802e9038",
  1044 => x"b9d80881",
  1045 => x"ff321281",
  1046 => x"05b9c40c",
  1047 => x"a1900471",
  1048 => x"b9d80831",
  1049 => x"b9c40ca1",
  1050 => x"9004b3e8",
  1051 => x"08ff05b3",
  1052 => x"e80cb3e8",
  1053 => x"08ff2e09",
  1054 => x"81069538",
  1055 => x"b3ec0880",
  1056 => x"2e8a3887",
  1057 => x"0bb3e408",
  1058 => x"31b3e40c",
  1059 => x"70b3ec0c",
  1060 => x"738a2a70",
  1061 => x"81065151",
  1062 => x"70802e92",
  1063 => x"38b3e008",
  1064 => x"51ff7125",
  1065 => x"893870e4",
  1066 => x"0cff0bb3",
  1067 => x"e00c800b",
  1068 => x"b9d00ca4",
  1069 => x"812da488",
  1070 => x"2d029005",
  1071 => x"0d0402fc",
  1072 => x"050db3e0",
  1073 => x"08517080",
  1074 => x"24fc3872",
  1075 => x"b3e00c02",
  1076 => x"84050d04",
  1077 => x"02fc050d",
  1078 => x"a48e2d81",
  1079 => x"0bb9d00c",
  1080 => x"a4882db9",
  1081 => x"d0085170",
  1082 => x"fa380284",
  1083 => x"050d0402",
  1084 => x"fc050db9",
  1085 => x"9c519ec7",
  1086 => x"2d9f9e51",
  1087 => x"a3fd2da3",
  1088 => x"a72d81f4",
  1089 => x"51a1be2d",
  1090 => x"0284050d",
  1091 => x"0402f405",
  1092 => x"0da38f04",
  1093 => x"b4bc0881",
  1094 => x"f02e0981",
  1095 => x"06893881",
  1096 => x"0bb4b00c",
  1097 => x"a38f04b4",
  1098 => x"bc0881e0",
  1099 => x"2e098106",
  1100 => x"8938810b",
  1101 => x"b4b40ca3",
  1102 => x"8f04b4bc",
  1103 => x"0852b4b4",
  1104 => x"08802e88",
  1105 => x"38b4bc08",
  1106 => x"81800552",
  1107 => x"71842c72",
  1108 => x"8f065353",
  1109 => x"b4b00880",
  1110 => x"2e993872",
  1111 => x"8429b3f0",
  1112 => x"05721381",
  1113 => x"712b7009",
  1114 => x"73080673",
  1115 => x"0c515353",
  1116 => x"a3850472",
  1117 => x"8429b3f0",
  1118 => x"05721383",
  1119 => x"712b7208",
  1120 => x"07720c53",
  1121 => x"53800bb4",
  1122 => x"b40c800b",
  1123 => x"b4b00cb9",
  1124 => x"9c519eda",
  1125 => x"2db4bc08",
  1126 => x"ff24fef8",
  1127 => x"38800bb4",
  1128 => x"bc0c028c",
  1129 => x"050d0402",
  1130 => x"f8050db3",
  1131 => x"f0528f51",
  1132 => x"80727084",
  1133 => x"05540cff",
  1134 => x"11517080",
  1135 => x"25f23802",
  1136 => x"88050d04",
  1137 => x"02f0050d",
  1138 => x"7551a48e",
  1139 => x"2d70822c",
  1140 => x"fc06b3f0",
  1141 => x"1172109e",
  1142 => x"06710870",
  1143 => x"722a7083",
  1144 => x"0682742b",
  1145 => x"70097406",
  1146 => x"760c5451",
  1147 => x"56575351",
  1148 => x"53a4882d",
  1149 => x"71b4bc0c",
  1150 => x"0290050d",
  1151 => x"0471980c",
  1152 => x"04ffb008",
  1153 => x"b4bc0c04",
  1154 => x"810bffb0",
  1155 => x"0c04800b",
  1156 => x"ffb00c04",
  1157 => x"02fc050d",
  1158 => x"800bb4b8",
  1159 => x"0c805184",
  1160 => x"e52d0284",
  1161 => x"050d0402",
  1162 => x"ec050d76",
  1163 => x"54805287",
  1164 => x"0b881580",
  1165 => x"f52d5653",
  1166 => x"74722483",
  1167 => x"38a05372",
  1168 => x"5182ee2d",
  1169 => x"81128b15",
  1170 => x"80f52d54",
  1171 => x"52727225",
  1172 => x"de380294",
  1173 => x"050d0402",
  1174 => x"f0050db9",
  1175 => x"e8085481",
  1176 => x"f72d800b",
  1177 => x"b9ec0c73",
  1178 => x"08802e81",
  1179 => x"8038820b",
  1180 => x"b4d00cb9",
  1181 => x"ec088f06",
  1182 => x"b4cc0c73",
  1183 => x"08527183",
  1184 => x"2e963871",
  1185 => x"83268938",
  1186 => x"71812eaf",
  1187 => x"38a5d804",
  1188 => x"71852e9f",
  1189 => x"38a5d804",
  1190 => x"881480f5",
  1191 => x"2d841508",
  1192 => x"b1985354",
  1193 => x"5285f32d",
  1194 => x"71842913",
  1195 => x"70085252",
  1196 => x"a5dc0473",
  1197 => x"51a4a72d",
  1198 => x"a5d804b9",
  1199 => x"e4088815",
  1200 => x"082c7081",
  1201 => x"06515271",
  1202 => x"802e8738",
  1203 => x"b19c51a5",
  1204 => x"d504b1a0",
  1205 => x"5185f32d",
  1206 => x"84140851",
  1207 => x"85f32db9",
  1208 => x"ec088105",
  1209 => x"b9ec0c8c",
  1210 => x"1454a4e7",
  1211 => x"04029005",
  1212 => x"0d0471b9",
  1213 => x"e80ca4d7",
  1214 => x"2db9ec08",
  1215 => x"ff05b9f0",
  1216 => x"0c0402ec",
  1217 => x"050db9e8",
  1218 => x"085580f8",
  1219 => x"51a3c42d",
  1220 => x"b4bc0881",
  1221 => x"2a708106",
  1222 => x"5152719b",
  1223 => x"388751a3",
  1224 => x"c42db4bc",
  1225 => x"08812a70",
  1226 => x"81065152",
  1227 => x"71802eb1",
  1228 => x"38a6b704",
  1229 => x"a28d2d87",
  1230 => x"51a3c42d",
  1231 => x"b4bc08f4",
  1232 => x"38a6c704",
  1233 => x"a28d2d80",
  1234 => x"f851a3c4",
  1235 => x"2db4bc08",
  1236 => x"f338b4b8",
  1237 => x"08813270",
  1238 => x"b4b80c70",
  1239 => x"525284e5",
  1240 => x"2db4b808",
  1241 => x"a23880da",
  1242 => x"51a3c42d",
  1243 => x"81f551a3",
  1244 => x"c42d81f2",
  1245 => x"51a3c42d",
  1246 => x"81eb51a3",
  1247 => x"c42d81f4",
  1248 => x"51a3c42d",
  1249 => x"aacb0481",
  1250 => x"f551a3c4",
  1251 => x"2db4bc08",
  1252 => x"812a7081",
  1253 => x"06515271",
  1254 => x"802e8f38",
  1255 => x"b9f00852",
  1256 => x"71802e86",
  1257 => x"38ff12b9",
  1258 => x"f00c81f2",
  1259 => x"51a3c42d",
  1260 => x"b4bc0881",
  1261 => x"2a708106",
  1262 => x"51527180",
  1263 => x"2e9538b9",
  1264 => x"ec08ff05",
  1265 => x"b9f00854",
  1266 => x"52727225",
  1267 => x"86388113",
  1268 => x"b9f00cb9",
  1269 => x"f0087053",
  1270 => x"5473802e",
  1271 => x"8a388c15",
  1272 => x"ff155555",
  1273 => x"a7d90482",
  1274 => x"0bb4d00c",
  1275 => x"718f06b4",
  1276 => x"cc0c81eb",
  1277 => x"51a3c42d",
  1278 => x"b4bc0881",
  1279 => x"2a708106",
  1280 => x"51527180",
  1281 => x"2ead3874",
  1282 => x"08852e09",
  1283 => x"8106a438",
  1284 => x"881580f5",
  1285 => x"2dff0552",
  1286 => x"71881681",
  1287 => x"b72d7198",
  1288 => x"2b527180",
  1289 => x"25883880",
  1290 => x"0b881681",
  1291 => x"b72d7451",
  1292 => x"a4a72d81",
  1293 => x"f451a3c4",
  1294 => x"2db4bc08",
  1295 => x"812a7081",
  1296 => x"06515271",
  1297 => x"802eb338",
  1298 => x"7408852e",
  1299 => x"098106aa",
  1300 => x"38881580",
  1301 => x"f52d8105",
  1302 => x"52718816",
  1303 => x"81b72d71",
  1304 => x"81ff068b",
  1305 => x"1680f52d",
  1306 => x"54527272",
  1307 => x"27873872",
  1308 => x"881681b7",
  1309 => x"2d7451a4",
  1310 => x"a72d80da",
  1311 => x"51a3c42d",
  1312 => x"b4bc0881",
  1313 => x"2a708106",
  1314 => x"51527180",
  1315 => x"2e80fb38",
  1316 => x"b9e808b9",
  1317 => x"f0085553",
  1318 => x"73802e8a",
  1319 => x"388c13ff",
  1320 => x"155553a9",
  1321 => x"98047208",
  1322 => x"5271822e",
  1323 => x"a6387182",
  1324 => x"26893871",
  1325 => x"812ea538",
  1326 => x"aa8a0471",
  1327 => x"832ead38",
  1328 => x"71842e09",
  1329 => x"810680c2",
  1330 => x"38881308",
  1331 => x"51a5f22d",
  1332 => x"aa8a0488",
  1333 => x"13085271",
  1334 => x"2daa8a04",
  1335 => x"810b8814",
  1336 => x"082bb9e4",
  1337 => x"0832b9e4",
  1338 => x"0caa8704",
  1339 => x"881380f5",
  1340 => x"2d81058b",
  1341 => x"1480f52d",
  1342 => x"53547174",
  1343 => x"24833880",
  1344 => x"54738814",
  1345 => x"81b72da4",
  1346 => x"d72d8054",
  1347 => x"800bb4d0",
  1348 => x"0c738f06",
  1349 => x"b4cc0ca0",
  1350 => x"5273b9f0",
  1351 => x"082e0981",
  1352 => x"069838b9",
  1353 => x"ec08ff05",
  1354 => x"74327009",
  1355 => x"81057072",
  1356 => x"079f2a91",
  1357 => x"71315151",
  1358 => x"53537151",
  1359 => x"82ee2d81",
  1360 => x"14548e74",
  1361 => x"25c638b4",
  1362 => x"b8085271",
  1363 => x"b4bc0c02",
  1364 => x"94050d04",
  1365 => x"00ffffff",
  1366 => x"ff00ffff",
  1367 => x"ffff00ff",
  1368 => x"ffffff00",
  1369 => x"52657365",
  1370 => x"74000000",
  1371 => x"4f707469",
  1372 => x"6f6e7320",
  1373 => x"10000000",
  1374 => x"536f756e",
  1375 => x"64201000",
  1376 => x"54757262",
  1377 => x"6f202831",
  1378 => x"302e3734",
  1379 => x"4d487a29",
  1380 => x"00000000",
  1381 => x"4d6f7573",
  1382 => x"6520656d",
  1383 => x"756c6174",
  1384 => x"696f6e00",
  1385 => x"45786974",
  1386 => x"00000000",
  1387 => x"4d617374",
  1388 => x"65720000",
  1389 => x"4f504c4c",
  1390 => x"00000000",
  1391 => x"53434300",
  1392 => x"50534700",
  1393 => x"4261636b",
  1394 => x"00000000",
  1395 => x"5363616e",
  1396 => x"6c696e65",
  1397 => x"73000000",
  1398 => x"53442043",
  1399 => x"61726400",
  1400 => x"4a617061",
  1401 => x"6e657365",
  1402 => x"206b6579",
  1403 => x"626f6172",
  1404 => x"64206c61",
  1405 => x"796f7574",
  1406 => x"00000000",
  1407 => x"32303438",
  1408 => x"4c422052",
  1409 => x"414d0000",
  1410 => x"34303936",
  1411 => x"4b422052",
  1412 => x"414d0000",
  1413 => x"536c323a",
  1414 => x"204e6f6e",
  1415 => x"65000000",
  1416 => x"536c323a",
  1417 => x"20455345",
  1418 => x"2d534343",
  1419 => x"20314d42",
  1420 => x"2f534343",
  1421 => x"2d490000",
  1422 => x"536c323a",
  1423 => x"20455345",
  1424 => x"2d52414d",
  1425 => x"20314d42",
  1426 => x"2f415343",
  1427 => x"49493800",
  1428 => x"536c323a",
  1429 => x"20455345",
  1430 => x"2d52414d",
  1431 => x"20314d42",
  1432 => x"2f415343",
  1433 => x"49493136",
  1434 => x"00000000",
  1435 => x"536c313a",
  1436 => x"204e6f6e",
  1437 => x"65000000",
  1438 => x"536c313a",
  1439 => x"20455345",
  1440 => x"2d534343",
  1441 => x"20314d42",
  1442 => x"2f534343",
  1443 => x"2d490000",
  1444 => x"536c313a",
  1445 => x"204d6567",
  1446 => x"6152414d",
  1447 => x"00000000",
  1448 => x"56474120",
  1449 => x"2d203331",
  1450 => x"4b487a2c",
  1451 => x"20363048",
  1452 => x"7a000000",
  1453 => x"56474120",
  1454 => x"2d203331",
  1455 => x"4b487a2c",
  1456 => x"20353048",
  1457 => x"7a000000",
  1458 => x"5456202d",
  1459 => x"20343830",
  1460 => x"692c2036",
  1461 => x"30487a00",
  1462 => x"496e6974",
  1463 => x"69616c69",
  1464 => x"7a696e67",
  1465 => x"20534420",
  1466 => x"63617264",
  1467 => x"0a000000",
  1468 => x"53444843",
  1469 => x"20636172",
  1470 => x"64206465",
  1471 => x"74656374",
  1472 => x"65642062",
  1473 => x"7574206e",
  1474 => x"6f740a73",
  1475 => x"7570706f",
  1476 => x"72746564",
  1477 => x"3b206469",
  1478 => x"7361626c",
  1479 => x"696e6720",
  1480 => x"53442063",
  1481 => x"6172640a",
  1482 => x"10204f4b",
  1483 => x"0a000000",
  1484 => x"46617433",
  1485 => x"32206669",
  1486 => x"6c657379",
  1487 => x"7374656d",
  1488 => x"20646574",
  1489 => x"65637465",
  1490 => x"64206275",
  1491 => x"740a6e6f",
  1492 => x"74207375",
  1493 => x"70706f72",
  1494 => x"7465643b",
  1495 => x"20646973",
  1496 => x"61626c69",
  1497 => x"6e672053",
  1498 => x"44206361",
  1499 => x"72640a10",
  1500 => x"204f4b0a",
  1501 => x"00000000",
  1502 => x"54727969",
  1503 => x"6e67204d",
  1504 => x"53583342",
  1505 => x"494f532e",
  1506 => x"5359532e",
  1507 => x"2e2e0a00",
  1508 => x"4d535833",
  1509 => x"42494f53",
  1510 => x"53595300",
  1511 => x"54727969",
  1512 => x"6e672042",
  1513 => x"494f535f",
  1514 => x"4d32502e",
  1515 => x"524f4d2e",
  1516 => x"2e2e0a00",
  1517 => x"42494f53",
  1518 => x"5f4d3250",
  1519 => x"524f4d00",
  1520 => x"4f70656e",
  1521 => x"65642042",
  1522 => x"494f532c",
  1523 => x"206c6f61",
  1524 => x"64696e67",
  1525 => x"2e2e2e0a",
  1526 => x"00000000",
  1527 => x"52656164",
  1528 => x"20626c6f",
  1529 => x"636b2066",
  1530 => x"61696c65",
  1531 => x"640a0000",
  1532 => x"4c6f6164",
  1533 => x"696e6720",
  1534 => x"42494f53",
  1535 => x"20666169",
  1536 => x"6c65640a",
  1537 => x"00000000",
  1538 => x"52656164",
  1539 => x"206f6620",
  1540 => x"4d425220",
  1541 => x"6661696c",
  1542 => x"65640a00",
  1543 => x"46415431",
  1544 => x"36202020",
  1545 => x"00000000",
  1546 => x"46415433",
  1547 => x"32202020",
  1548 => x"00000000",
  1549 => x"4e6f2070",
  1550 => x"61727469",
  1551 => x"74696f6e",
  1552 => x"20736967",
  1553 => x"0a000000",
  1554 => x"42616420",
  1555 => x"70617274",
  1556 => x"0a000000",
  1557 => x"53444843",
  1558 => x"20657272",
  1559 => x"6f72210a",
  1560 => x"00000000",
  1561 => x"53442069",
  1562 => x"6e69742e",
  1563 => x"2e2e0a00",
  1564 => x"53442063",
  1565 => x"61726420",
  1566 => x"72657365",
  1567 => x"74206661",
  1568 => x"696c6564",
  1569 => x"210a0000",
  1570 => x"52656164",
  1571 => x"20666169",
  1572 => x"6c65640a",
  1573 => x"00000000",
  1574 => x"16200000",
  1575 => x"14200000",
  1576 => x"15200000",
  1577 => x"00000002",
  1578 => x"00000002",
  1579 => x"00001564",
  1580 => x"00000540",
  1581 => x"00000004",
  1582 => x"0000156c",
  1583 => x"00001944",
  1584 => x"00000004",
  1585 => x"00001578",
  1586 => x"000018fc",
  1587 => x"00000001",
  1588 => x"00001580",
  1589 => x"00000007",
  1590 => x"00000001",
  1591 => x"00001594",
  1592 => x"0000000a",
  1593 => x"00000002",
  1594 => x"000015a4",
  1595 => x"00001214",
  1596 => x"00000000",
  1597 => x"00000000",
  1598 => x"00000000",
  1599 => x"00000005",
  1600 => x"000015ac",
  1601 => x"00000007",
  1602 => x"00000005",
  1603 => x"000015b4",
  1604 => x"00000007",
  1605 => x"00000005",
  1606 => x"000015bc",
  1607 => x"00000007",
  1608 => x"00000005",
  1609 => x"000015c0",
  1610 => x"00000007",
  1611 => x"00000004",
  1612 => x"000015c4",
  1613 => x"000018a8",
  1614 => x"00000000",
  1615 => x"00000000",
  1616 => x"00000000",
  1617 => x"00000003",
  1618 => x"000019d4",
  1619 => x"00000003",
  1620 => x"00000001",
  1621 => x"000015cc",
  1622 => x"0000000b",
  1623 => x"00000001",
  1624 => x"000015d8",
  1625 => x"00000002",
  1626 => x"00000003",
  1627 => x"000019c8",
  1628 => x"00000003",
  1629 => x"00000003",
  1630 => x"000019b8",
  1631 => x"00000004",
  1632 => x"00000001",
  1633 => x"000015e0",
  1634 => x"00000006",
  1635 => x"00000003",
  1636 => x"000019b0",
  1637 => x"00000002",
  1638 => x"00000004",
  1639 => x"000015c4",
  1640 => x"000018a8",
  1641 => x"00000000",
  1642 => x"00000000",
  1643 => x"00000000",
  1644 => x"000015fc",
  1645 => x"00001608",
  1646 => x"00001614",
  1647 => x"00001620",
  1648 => x"00001638",
  1649 => x"00001650",
  1650 => x"0000166c",
  1651 => x"00001678",
  1652 => x"00001690",
  1653 => x"000016a0",
  1654 => x"000016b4",
  1655 => x"000016c8",
  1656 => x"ffffffff",
  1657 => x"00000003",
  1658 => x"00000000",
  1659 => x"00000000",
  1660 => x"00000000",
  1661 => x"00000000",
  1662 => x"00000000",
  1663 => x"00000000",
  1664 => x"00000000",
  1665 => x"00000000",
  1666 => x"00000000",
  1667 => x"00000000",
  1668 => x"00000000",
  1669 => x"00000000",
  1670 => x"00000000",
  1671 => x"00000000",
  1672 => x"00000000",
  1673 => x"00000000",
  1674 => x"00000000",
  1675 => x"00000000",
  1676 => x"00000000",
  1677 => x"00000000",
  1678 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

