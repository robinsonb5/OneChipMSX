-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b0bb2",
     9 => x"e8080b0b",
    10 => x"0bb2ec08",
    11 => x"0b0b0bb2",
    12 => x"f0080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"b2f00c0b",
    16 => x"0b0bb2ec",
    17 => x"0c0b0b0b",
    18 => x"b2e80c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0ba394",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"b2e870b9",
    57 => x"c4278b38",
    58 => x"80717084",
    59 => x"05530c81",
    60 => x"e2048c51",
    61 => x"81f70402",
    62 => x"dc050db9",
    63 => x"0bd00c81",
    64 => x"0bd40c84",
    65 => x"0bd40ca3",
    66 => x"a45195bf",
    67 => x"2d92e02d",
    68 => x"b2e80880",
    69 => x"2e81a638",
    70 => x"a3bc5195",
    71 => x"bf2d849f",
    72 => x"2da3d452",
    73 => x"b4a0518b",
    74 => x"842db2e8",
    75 => x"0881ff06",
    76 => x"5372802e",
    77 => x"818138a3",
    78 => x"e05195bf",
    79 => x"2db4a408",
    80 => x"83ff0589",
    81 => x"2a538073",
    82 => x"2580f238",
    83 => x"7258ae51",
    84 => x"959d2db4",
    85 => x"b852b4a0",
    86 => x"518ddf2d",
    87 => x"b2e80881",
    88 => x"ff065372",
    89 => x"802eba38",
    90 => x"b4b85983",
    91 => x"fc577870",
    92 => x"84055a08",
    93 => x"70828029",
    94 => x"71317188",
    95 => x"2c7081ff",
    96 => x"0673902c",
    97 => x"7081ff06",
    98 => x"75982ad8",
    99 => x"0cd80c58",
   100 => x"d80c57d8",
   101 => x"0cfc1858",
   102 => x"53768025",
   103 => x"d13883a7",
   104 => x"04a3fc51",
   105 => x"95bf2db4",
   106 => x"a0518db2",
   107 => x"2dff1858",
   108 => x"77ff9b38",
   109 => x"83bd04a4",
   110 => x"905195bf",
   111 => x"2d800bd4",
   112 => x"0ca4a851",
   113 => x"95bf2d9e",
   114 => x"e82da296",
   115 => x"2d9f802d",
   116 => x"b2e80880",
   117 => x"2ef738b2",
   118 => x"e8085195",
   119 => x"9d2d83cd",
   120 => x"0402e805",
   121 => x"0d77797b",
   122 => x"58555580",
   123 => x"53727625",
   124 => x"a3387470",
   125 => x"81055680",
   126 => x"f52d7470",
   127 => x"81055680",
   128 => x"f52d5252",
   129 => x"71712e86",
   130 => x"38815184",
   131 => x"96048113",
   132 => x"5383ed04",
   133 => x"805170b2",
   134 => x"e80c0298",
   135 => x"050d0402",
   136 => x"d8050dff",
   137 => x"0bb8c00c",
   138 => x"800bb8d4",
   139 => x"0ca4c851",
   140 => x"95bf2db4",
   141 => x"b8528051",
   142 => x"93fa2db2",
   143 => x"e80854b2",
   144 => x"e8088c38",
   145 => x"a4d85195",
   146 => x"bf2d7355",
   147 => x"89f704a4",
   148 => x"ec5195bf",
   149 => x"2d805681",
   150 => x"0bb4ac0c",
   151 => x"8853a584",
   152 => x"52b4ee51",
   153 => x"83e12db2",
   154 => x"e808762e",
   155 => x"09810687",
   156 => x"38b2e808",
   157 => x"b4ac0c88",
   158 => x"53a59052",
   159 => x"b58a5183",
   160 => x"e12db2e8",
   161 => x"088738b2",
   162 => x"e808b4ac",
   163 => x"0cb4ac08",
   164 => x"52a59c51",
   165 => x"97c72db4",
   166 => x"ac08802e",
   167 => x"818738b7",
   168 => x"fe0b80f5",
   169 => x"2db7ff0b",
   170 => x"80f52d71",
   171 => x"982b7190",
   172 => x"2b07b880",
   173 => x"0b80f52d",
   174 => x"70882b72",
   175 => x"07b8810b",
   176 => x"80f52d71",
   177 => x"07b8b60b",
   178 => x"80f52db8",
   179 => x"b70b80f5",
   180 => x"2d71882b",
   181 => x"07535f54",
   182 => x"525a5657",
   183 => x"557381ab",
   184 => x"aa2e0981",
   185 => x"068d3875",
   186 => x"5196872d",
   187 => x"b2e80856",
   188 => x"86830473",
   189 => x"82d4d52e",
   190 => x"8a38a5b0",
   191 => x"5195bf2d",
   192 => x"87b80475",
   193 => x"52a5d051",
   194 => x"97c72db4",
   195 => x"b8527551",
   196 => x"93fa2db2",
   197 => x"e80855b2",
   198 => x"e808802e",
   199 => x"83d938a5",
   200 => x"e85195bf",
   201 => x"2da69051",
   202 => x"97c72d88",
   203 => x"53a59052",
   204 => x"b58a5183",
   205 => x"e12db2e8",
   206 => x"08893881",
   207 => x"0bb8d40c",
   208 => x"86de0488",
   209 => x"53a58452",
   210 => x"b4ee5183",
   211 => x"e12db2e8",
   212 => x"08802e8a",
   213 => x"38a6a851",
   214 => x"97c72d87",
   215 => x"b804b8b6",
   216 => x"0b80f52d",
   217 => x"547380d5",
   218 => x"2e098106",
   219 => x"80ca38b8",
   220 => x"b70b80f5",
   221 => x"2d547381",
   222 => x"aa2e0981",
   223 => x"06ba3880",
   224 => x"0bb4b80b",
   225 => x"80f52d56",
   226 => x"547481e9",
   227 => x"2e833881",
   228 => x"547481eb",
   229 => x"2e8c3880",
   230 => x"5573752e",
   231 => x"09810682",
   232 => x"d638b4c3",
   233 => x"0b80f52d",
   234 => x"59788d38",
   235 => x"b4c40b80",
   236 => x"f52d5473",
   237 => x"822e8638",
   238 => x"805589f7",
   239 => x"04b4c50b",
   240 => x"80f52d70",
   241 => x"b8dc0cff",
   242 => x"1170b8d0",
   243 => x"0c5452a6",
   244 => x"c85197c7",
   245 => x"2db4c60b",
   246 => x"80f52db4",
   247 => x"c70b80f5",
   248 => x"2d567605",
   249 => x"75828029",
   250 => x"0570b8c4",
   251 => x"0cb4c80b",
   252 => x"80f52d70",
   253 => x"b8bc0cb8",
   254 => x"d4085957",
   255 => x"5876802e",
   256 => x"81a53888",
   257 => x"53a59052",
   258 => x"b58a5183",
   259 => x"e12d7855",
   260 => x"b2e80881",
   261 => x"e238b8dc",
   262 => x"0870842b",
   263 => x"b8b80c70",
   264 => x"b8d80cb4",
   265 => x"dd0b80f5",
   266 => x"2db4dc0b",
   267 => x"80f52d71",
   268 => x"82802905",
   269 => x"b4de0b80",
   270 => x"f52d7084",
   271 => x"80802912",
   272 => x"b4df0b80",
   273 => x"f52d7081",
   274 => x"800a2912",
   275 => x"70b4b00c",
   276 => x"b8bc0871",
   277 => x"29b8c408",
   278 => x"0570b8e4",
   279 => x"0cb4e50b",
   280 => x"80f52db4",
   281 => x"e40b80f5",
   282 => x"2d718280",
   283 => x"2905b4e6",
   284 => x"0b80f52d",
   285 => x"70848080",
   286 => x"2912b4e7",
   287 => x"0b80f52d",
   288 => x"70982b81",
   289 => x"f00a0672",
   290 => x"0570b4b4",
   291 => x"0cfe117e",
   292 => x"297705b8",
   293 => x"cc0c5257",
   294 => x"52575d57",
   295 => x"51525f52",
   296 => x"5c575757",
   297 => x"89f504b4",
   298 => x"ca0b80f5",
   299 => x"2db4c90b",
   300 => x"80f52d71",
   301 => x"82802905",
   302 => x"70b8b80c",
   303 => x"70a02983",
   304 => x"ff057089",
   305 => x"2a70b8d8",
   306 => x"0cb4cf0b",
   307 => x"80f52db4",
   308 => x"ce0b80f5",
   309 => x"2d718280",
   310 => x"290570b4",
   311 => x"b00c7b71",
   312 => x"291e70b8",
   313 => x"cc0c7db4",
   314 => x"b40c7305",
   315 => x"b8e40c55",
   316 => x"5e515155",
   317 => x"55815574",
   318 => x"b2e80c02",
   319 => x"a8050d04",
   320 => x"02ec050d",
   321 => x"7670872c",
   322 => x"7180ff06",
   323 => x"575553b8",
   324 => x"d4088a38",
   325 => x"72882c73",
   326 => x"81ff0656",
   327 => x"5473b8c0",
   328 => x"082ea638",
   329 => x"b8c40814",
   330 => x"52a6ec51",
   331 => x"97c72db4",
   332 => x"b852b8c4",
   333 => x"08145193",
   334 => x"fa2db2e8",
   335 => x"0853b2e8",
   336 => x"08802eb7",
   337 => x"3873b8c0",
   338 => x"0cb8d408",
   339 => x"802e9838",
   340 => x"748429b4",
   341 => x"b8057008",
   342 => x"52539687",
   343 => x"2db2e808",
   344 => x"f00a0655",
   345 => x"8af90474",
   346 => x"10b4b805",
   347 => x"7080e02d",
   348 => x"525396b7",
   349 => x"2db2e808",
   350 => x"55745372",
   351 => x"b2e80c02",
   352 => x"94050d04",
   353 => x"02c8050d",
   354 => x"7f615f5c",
   355 => x"8057ff0b",
   356 => x"b8c00cb4",
   357 => x"b408b8cc",
   358 => x"085758b8",
   359 => x"d408772e",
   360 => x"8a38b8dc",
   361 => x"08842b59",
   362 => x"8bb104b8",
   363 => x"d808842b",
   364 => x"59805a79",
   365 => x"792781b6",
   366 => x"38798f06",
   367 => x"a0185854",
   368 => x"73973875",
   369 => x"52a78c51",
   370 => x"97c72db4",
   371 => x"b8527551",
   372 => x"81165693",
   373 => x"fa2db4b8",
   374 => x"57807780",
   375 => x"f52d5654",
   376 => x"74742e83",
   377 => x"38815474",
   378 => x"81e52e80",
   379 => x"fb388170",
   380 => x"7506555d",
   381 => x"73802e80",
   382 => x"ef388b17",
   383 => x"80f52d98",
   384 => x"065b7a80",
   385 => x"e3387651",
   386 => x"95bf2d8b",
   387 => x"537d5276",
   388 => x"5183e12d",
   389 => x"b2e80880",
   390 => x"cf389c17",
   391 => x"08519687",
   392 => x"2db2e808",
   393 => x"841d0c9a",
   394 => x"1780e02d",
   395 => x"5196b72d",
   396 => x"b2e808b2",
   397 => x"e808881e",
   398 => x"0cb2e808",
   399 => x"5555b8d4",
   400 => x"08802e98",
   401 => x"38941780",
   402 => x"e02d5196",
   403 => x"b72db2e8",
   404 => x"08902b83",
   405 => x"fff00a06",
   406 => x"70165154",
   407 => x"73881d0c",
   408 => x"7a7c0c7c",
   409 => x"548da904",
   410 => x"811a5a8b",
   411 => x"b304b8d4",
   412 => x"08802eb3",
   413 => x"3877518a",
   414 => x"802db2e8",
   415 => x"08b2e808",
   416 => x"53a7ac52",
   417 => x"5897c72d",
   418 => x"7780ffff",
   419 => x"fff80654",
   420 => x"7380ffff",
   421 => x"fff82e8f",
   422 => x"38fe18b8",
   423 => x"dc0829b8",
   424 => x"e4080556",
   425 => x"8bb10480",
   426 => x"5473b2e8",
   427 => x"0c02b805",
   428 => x"0d0402f4",
   429 => x"050d7470",
   430 => x"08810571",
   431 => x"0c7008b8",
   432 => x"d0080653",
   433 => x"53718e38",
   434 => x"88130851",
   435 => x"8a802db2",
   436 => x"e8088814",
   437 => x"0c810bb2",
   438 => x"e80c028c",
   439 => x"050d0402",
   440 => x"f0050d75",
   441 => x"881108fe",
   442 => x"05b8dc08",
   443 => x"29b8e408",
   444 => x"117208b8",
   445 => x"d0080605",
   446 => x"79555354",
   447 => x"5493fa2d",
   448 => x"b2e80853",
   449 => x"b2e80880",
   450 => x"2e833881",
   451 => x"5372b2e8",
   452 => x"0c029005",
   453 => x"0d0402f4",
   454 => x"050dd452",
   455 => x"81ff720c",
   456 => x"71085381",
   457 => x"ff720c72",
   458 => x"882b83fe",
   459 => x"80067208",
   460 => x"7081ff06",
   461 => x"51525381",
   462 => x"ff720c72",
   463 => x"7107882b",
   464 => x"72087081",
   465 => x"ff065152",
   466 => x"5381ff72",
   467 => x"0c727107",
   468 => x"882b7208",
   469 => x"7081ff06",
   470 => x"7207b2e8",
   471 => x"0c525302",
   472 => x"8c050d04",
   473 => x"02f4050d",
   474 => x"74767181",
   475 => x"ff06d40c",
   476 => x"5353b8e8",
   477 => x"08853871",
   478 => x"892b5271",
   479 => x"982ad40c",
   480 => x"71902a70",
   481 => x"81ff06d4",
   482 => x"0c517188",
   483 => x"2a7081ff",
   484 => x"06d40c51",
   485 => x"7181ff06",
   486 => x"d40c7290",
   487 => x"2a7081ff",
   488 => x"06d40c51",
   489 => x"d4087081",
   490 => x"ff065151",
   491 => x"82b8bf52",
   492 => x"7081ff2e",
   493 => x"09810694",
   494 => x"3881ff0b",
   495 => x"d40cd408",
   496 => x"7081ff06",
   497 => x"ff145451",
   498 => x"5171e538",
   499 => x"70b2e80c",
   500 => x"028c050d",
   501 => x"0402fc05",
   502 => x"0d81c751",
   503 => x"81ff0bd4",
   504 => x"0cff1151",
   505 => x"708025f4",
   506 => x"38028405",
   507 => x"0d0402f0",
   508 => x"050d8fd5",
   509 => x"2d819c9f",
   510 => x"53805287",
   511 => x"fc80f751",
   512 => x"8ee42db2",
   513 => x"e80854b2",
   514 => x"e808812e",
   515 => x"098106a3",
   516 => x"3881ff0b",
   517 => x"d40c820a",
   518 => x"52849c80",
   519 => x"e9518ee4",
   520 => x"2db2e808",
   521 => x"8b3881ff",
   522 => x"0bd40c73",
   523 => x"5390b904",
   524 => x"8fd52dff",
   525 => x"135372c1",
   526 => x"3872b2e8",
   527 => x"0c029005",
   528 => x"0d0402f4",
   529 => x"050d81ff",
   530 => x"0bd40ca7",
   531 => x"c45195bf",
   532 => x"2d935380",
   533 => x"5287fc80",
   534 => x"c1518ee4",
   535 => x"2db2e808",
   536 => x"8b3881ff",
   537 => x"0bd40c81",
   538 => x"5390f504",
   539 => x"8fd52dff",
   540 => x"135372df",
   541 => x"3872b2e8",
   542 => x"0c028c05",
   543 => x"0d0402f0",
   544 => x"050d8fd5",
   545 => x"2d83aa52",
   546 => x"849c80c8",
   547 => x"518ee42d",
   548 => x"b2e808b2",
   549 => x"e80853a7",
   550 => x"d0525397",
   551 => x"c72d7281",
   552 => x"2e098106",
   553 => x"9c388e96",
   554 => x"2db2e808",
   555 => x"83ffff06",
   556 => x"537283aa",
   557 => x"2ea138b2",
   558 => x"e80852a7",
   559 => x"e85197c7",
   560 => x"2d90c22d",
   561 => x"91d20481",
   562 => x"5492d704",
   563 => x"a8805197",
   564 => x"c72d8054",
   565 => x"92d70481",
   566 => x"ff0bd40c",
   567 => x"b1538fee",
   568 => x"2db2e808",
   569 => x"802e80e0",
   570 => x"38805287",
   571 => x"fc80fa51",
   572 => x"8ee42db2",
   573 => x"e80880c6",
   574 => x"38b2e808",
   575 => x"52a89c51",
   576 => x"97c72d81",
   577 => x"ff0bd40c",
   578 => x"d4087081",
   579 => x"ff067054",
   580 => x"a8a85351",
   581 => x"5397c72d",
   582 => x"81ff0bd4",
   583 => x"0c81ff0b",
   584 => x"d40c81ff",
   585 => x"0bd40c81",
   586 => x"ff0bd40c",
   587 => x"72862a70",
   588 => x"81067056",
   589 => x"51537280",
   590 => x"2e9d3891",
   591 => x"c704b2e8",
   592 => x"0852a89c",
   593 => x"5197c72d",
   594 => x"72822efe",
   595 => x"ff38ff13",
   596 => x"5372ff8a",
   597 => x"38725473",
   598 => x"b2e80c02",
   599 => x"90050d04",
   600 => x"02f4050d",
   601 => x"810bb8e8",
   602 => x"0cd00870",
   603 => x"8f2a7081",
   604 => x"06515153",
   605 => x"72f33872",
   606 => x"d00c8fd5",
   607 => x"2da8b851",
   608 => x"95bf2dd0",
   609 => x"08708f2a",
   610 => x"70810651",
   611 => x"515372f3",
   612 => x"38810bd0",
   613 => x"0c875380",
   614 => x"5284d480",
   615 => x"c0518ee4",
   616 => x"2db2e808",
   617 => x"812e9438",
   618 => x"72822e09",
   619 => x"81068638",
   620 => x"805393eb",
   621 => x"04ff1353",
   622 => x"72dd3890",
   623 => x"fe2db2e8",
   624 => x"08b8e80c",
   625 => x"815287fc",
   626 => x"80d0518e",
   627 => x"e42d81ff",
   628 => x"0bd40cd0",
   629 => x"08708f2a",
   630 => x"70810651",
   631 => x"515372f3",
   632 => x"3872d00c",
   633 => x"81ff0bd4",
   634 => x"0c815372",
   635 => x"b2e80c02",
   636 => x"8c050d04",
   637 => x"800bb2e8",
   638 => x"0c0402e0",
   639 => x"050d797b",
   640 => x"57578058",
   641 => x"81ff0bd4",
   642 => x"0cd00870",
   643 => x"8f2a7081",
   644 => x"06515154",
   645 => x"73f33882",
   646 => x"810bd00c",
   647 => x"81ff0bd4",
   648 => x"0c765287",
   649 => x"fc80d151",
   650 => x"8ee42d80",
   651 => x"dbc6df55",
   652 => x"b2e80880",
   653 => x"2e9038b2",
   654 => x"e8085376",
   655 => x"52a8c451",
   656 => x"97c72d95",
   657 => x"940481ff",
   658 => x"0bd40cd4",
   659 => x"087081ff",
   660 => x"06515473",
   661 => x"81fe2e09",
   662 => x"81069d38",
   663 => x"80ff548e",
   664 => x"962db2e8",
   665 => x"08767084",
   666 => x"05580cff",
   667 => x"14547380",
   668 => x"25ed3881",
   669 => x"5894fe04",
   670 => x"ff155574",
   671 => x"c93881ff",
   672 => x"0bd40cd0",
   673 => x"08708f2a",
   674 => x"70810651",
   675 => x"515473f3",
   676 => x"3873d00c",
   677 => x"77b2e80c",
   678 => x"02a0050d",
   679 => x"0402f805",
   680 => x"0d7352c0",
   681 => x"0870882a",
   682 => x"70810651",
   683 => x"51517080",
   684 => x"2ef13871",
   685 => x"c00c71b2",
   686 => x"e80c0288",
   687 => x"050d0402",
   688 => x"e8050d80",
   689 => x"78575575",
   690 => x"70840557",
   691 => x"08538054",
   692 => x"72982a73",
   693 => x"882b5452",
   694 => x"71802ea2",
   695 => x"38c00870",
   696 => x"882a7081",
   697 => x"06515151",
   698 => x"70802ef1",
   699 => x"3871c00c",
   700 => x"81158115",
   701 => x"55558374",
   702 => x"25d63871",
   703 => x"ca3874b2",
   704 => x"e80c0298",
   705 => x"050d0402",
   706 => x"f4050d74",
   707 => x"70882a83",
   708 => x"fe800670",
   709 => x"72982a07",
   710 => x"72882b87",
   711 => x"fc808006",
   712 => x"73982b81",
   713 => x"f00a0671",
   714 => x"730707b2",
   715 => x"e80c5651",
   716 => x"5351028c",
   717 => x"050d0402",
   718 => x"f8050d02",
   719 => x"8e0580f5",
   720 => x"2d74882b",
   721 => x"077083ff",
   722 => x"ff06b2e8",
   723 => x"0c510288",
   724 => x"050d0402",
   725 => x"f8050d73",
   726 => x"70902b71",
   727 => x"902a07b2",
   728 => x"e80c5202",
   729 => x"88050d04",
   730 => x"02ec050d",
   731 => x"76538055",
   732 => x"7275258b",
   733 => x"38ad5195",
   734 => x"9d2d7209",
   735 => x"81055372",
   736 => x"802eb538",
   737 => x"8754729c",
   738 => x"2a73842b",
   739 => x"54527180",
   740 => x"2e833881",
   741 => x"55897225",
   742 => x"8738b712",
   743 => x"5297a304",
   744 => x"b0125274",
   745 => x"802e8638",
   746 => x"7151959d",
   747 => x"2dff1454",
   748 => x"738025d2",
   749 => x"3897bd04",
   750 => x"b051959d",
   751 => x"2d800bb2",
   752 => x"e80c0294",
   753 => x"050d0402",
   754 => x"c0050d02",
   755 => x"80c40557",
   756 => x"80707870",
   757 => x"84055a08",
   758 => x"72415f5d",
   759 => x"587c7084",
   760 => x"055e085a",
   761 => x"805b7998",
   762 => x"2a7a882b",
   763 => x"5b567586",
   764 => x"38775f99",
   765 => x"bf047d80",
   766 => x"2e81a238",
   767 => x"805e7580",
   768 => x"e42e8a38",
   769 => x"7580f82e",
   770 => x"09810689",
   771 => x"38768418",
   772 => x"71085e58",
   773 => x"547580e4",
   774 => x"2e9f3875",
   775 => x"80e4268a",
   776 => x"387580e3",
   777 => x"2ebe3898",
   778 => x"ef047580",
   779 => x"f32ea338",
   780 => x"7580f82e",
   781 => x"893898ef",
   782 => x"048a5398",
   783 => x"c0049053",
   784 => x"b3c8527b",
   785 => x"5196e82d",
   786 => x"b2e808b3",
   787 => x"c85a5598",
   788 => x"ff047684",
   789 => x"18710870",
   790 => x"545b5854",
   791 => x"95bf2d80",
   792 => x"5598ff04",
   793 => x"76841871",
   794 => x"08585854",
   795 => x"99aa04a5",
   796 => x"51959d2d",
   797 => x"7551959d",
   798 => x"2d821858",
   799 => x"99b20474",
   800 => x"ff165654",
   801 => x"807425aa",
   802 => x"38787081",
   803 => x"055a80f5",
   804 => x"2d705256",
   805 => x"959d2d81",
   806 => x"185898ff",
   807 => x"0475a52e",
   808 => x"09810686",
   809 => x"38815e99",
   810 => x"b2047551",
   811 => x"959d2d81",
   812 => x"1858811b",
   813 => x"5b837b25",
   814 => x"feac3875",
   815 => x"fe9f387e",
   816 => x"b2e80c02",
   817 => x"80c0050d",
   818 => x"0402ec05",
   819 => x"0d765574",
   820 => x"80f52d51",
   821 => x"70802e81",
   822 => x"f238b48c",
   823 => x"08708280",
   824 => x"8029a8e4",
   825 => x"0805b488",
   826 => x"08115152",
   827 => x"52718f24",
   828 => x"de387470",
   829 => x"81055680",
   830 => x"f52d5271",
   831 => x"802e81cb",
   832 => x"3871882e",
   833 => x"0981069c",
   834 => x"38800bb4",
   835 => x"880825b8",
   836 => x"38ff1151",
   837 => x"a07181b7",
   838 => x"2db48808",
   839 => x"ff05b488",
   840 => x"0c9af004",
   841 => x"718a2e09",
   842 => x"81069d38",
   843 => x"b48c0881",
   844 => x"05b48c0c",
   845 => x"800bb488",
   846 => x"0cb48c08",
   847 => x"82808029",
   848 => x"a8e40805",
   849 => x"519af004",
   850 => x"71717081",
   851 => x"055381b7",
   852 => x"2db48808",
   853 => x"8105b488",
   854 => x"0cb48808",
   855 => x"a02e0981",
   856 => x"068e3880",
   857 => x"0bb4880c",
   858 => x"b48c0881",
   859 => x"05b48c0c",
   860 => x"8f0bb48c",
   861 => x"082580c7",
   862 => x"38a8e408",
   863 => x"82808011",
   864 => x"71535553",
   865 => x"81ff5273",
   866 => x"70840555",
   867 => x"08717084",
   868 => x"05530cff",
   869 => x"12527180",
   870 => x"25ed3888",
   871 => x"8013518f",
   872 => x"52807170",
   873 => x"8405530c",
   874 => x"ff125271",
   875 => x"8025f238",
   876 => x"800bb488",
   877 => x"0c8f0bb4",
   878 => x"8c0c9e80",
   879 => x"8013518f",
   880 => x"0bb48c08",
   881 => x"25feab38",
   882 => x"99cf0402",
   883 => x"94050d04",
   884 => x"02f4050d",
   885 => x"02930580",
   886 => x"f52d028c",
   887 => x"0581b72d",
   888 => x"80028405",
   889 => x"890581b7",
   890 => x"2d028c05",
   891 => x"fc055199",
   892 => x"c92d810b",
   893 => x"b2e80c02",
   894 => x"8c050d04",
   895 => x"02fc050d",
   896 => x"725199c9",
   897 => x"2d800bb2",
   898 => x"e80c0284",
   899 => x"050d0402",
   900 => x"f8050da8",
   901 => x"e408528f",
   902 => x"fc518072",
   903 => x"70840554",
   904 => x"0cfc1151",
   905 => x"708025f2",
   906 => x"38028805",
   907 => x"0d0402fc",
   908 => x"050d7251",
   909 => x"80710c80",
   910 => x"0b84120c",
   911 => x"800b8812",
   912 => x"0c800b8c",
   913 => x"120c0284",
   914 => x"050d0402",
   915 => x"f0050d75",
   916 => x"70088412",
   917 => x"08535353",
   918 => x"ff547171",
   919 => x"2e9b3884",
   920 => x"13087084",
   921 => x"29149311",
   922 => x"80f52d84",
   923 => x"16088111",
   924 => x"87068418",
   925 => x"0c525651",
   926 => x"5173b2e8",
   927 => x"0c029005",
   928 => x"0d0402f4",
   929 => x"050d7470",
   930 => x"08841208",
   931 => x"53535370",
   932 => x"72248f38",
   933 => x"72088414",
   934 => x"08717131",
   935 => x"5252529d",
   936 => x"af047208",
   937 => x"84140871",
   938 => x"71318805",
   939 => x"52525271",
   940 => x"b2e80c02",
   941 => x"8c050d04",
   942 => x"02f8050d",
   943 => x"a29c2da2",
   944 => x"8f2de008",
   945 => x"708b2a70",
   946 => x"81065152",
   947 => x"5270802e",
   948 => x"9d38b8f4",
   949 => x"08708429",
   950 => x"b9840573",
   951 => x"81ff0671",
   952 => x"0c5151b8",
   953 => x"f4088111",
   954 => x"8706b8f4",
   955 => x"0c51718a",
   956 => x"2a708106",
   957 => x"51517080",
   958 => x"2ea838b8",
   959 => x"fc08b980",
   960 => x"08525271",
   961 => x"712e9b38",
   962 => x"b8fc0870",
   963 => x"8429b9a4",
   964 => x"057008e0",
   965 => x"0c5151b8",
   966 => x"fc088111",
   967 => x"8706b8fc",
   968 => x"0c51a296",
   969 => x"2d028805",
   970 => x"0d0402f4",
   971 => x"050d7453",
   972 => x"8c130881",
   973 => x"11870688",
   974 => x"15085451",
   975 => x"5171712e",
   976 => x"ef38a29c",
   977 => x"2d8c1308",
   978 => x"70842914",
   979 => x"77b0120c",
   980 => x"51518c13",
   981 => x"08811187",
   982 => x"068c150c",
   983 => x"519db82d",
   984 => x"a2962d02",
   985 => x"8c050d04",
   986 => x"02fc050d",
   987 => x"b8f4519c",
   988 => x"ae2d9db8",
   989 => x"51a28b2d",
   990 => x"a1c32d02",
   991 => x"84050d04",
   992 => x"02e4050d",
   993 => x"8057a18e",
   994 => x"04b2e808",
   995 => x"81f02e09",
   996 => x"81068938",
   997 => x"810bb498",
   998 => x"0ca18e04",
   999 => x"b2e80881",
  1000 => x"e02e0981",
  1001 => x"06893881",
  1002 => x"0bb49c0c",
  1003 => x"a18e04b2",
  1004 => x"e80854b4",
  1005 => x"9c08802e",
  1006 => x"8838b2e8",
  1007 => x"08818005",
  1008 => x"54b49808",
  1009 => x"819c3883",
  1010 => x"0ba8e815",
  1011 => x"81b72d74",
  1012 => x"80ff24b1",
  1013 => x"38b49408",
  1014 => x"822a7081",
  1015 => x"06b49008",
  1016 => x"70872b81",
  1017 => x"80077811",
  1018 => x"822b5156",
  1019 => x"58515473",
  1020 => x"8b387581",
  1021 => x"80291570",
  1022 => x"822b5153",
  1023 => x"aae81308",
  1024 => x"537281b6",
  1025 => x"38800bb4",
  1026 => x"9c0c7480",
  1027 => x"d92e80c7",
  1028 => x"387480d9",
  1029 => x"248f3874",
  1030 => x"922ebc38",
  1031 => x"7480d82e",
  1032 => x"9338a189",
  1033 => x"047480f7",
  1034 => x"2ea03874",
  1035 => x"80fe2e8f",
  1036 => x"38a18904",
  1037 => x"b4940884",
  1038 => x"32b4940c",
  1039 => x"a0d204b4",
  1040 => x"94088132",
  1041 => x"b4940ca0",
  1042 => x"d204b494",
  1043 => x"088232b4",
  1044 => x"940c8157",
  1045 => x"a18904b4",
  1046 => x"90088107",
  1047 => x"b4900ca1",
  1048 => x"8904a8e8",
  1049 => x"1480f52d",
  1050 => x"81fe0653",
  1051 => x"72a8e815",
  1052 => x"81b72d74",
  1053 => x"922e8a38",
  1054 => x"7480d92e",
  1055 => x"09810689",
  1056 => x"38b49008",
  1057 => x"fe06b490",
  1058 => x"0c800bb4",
  1059 => x"980cb8f4",
  1060 => x"519ccb2d",
  1061 => x"b2e80855",
  1062 => x"b2e808ff",
  1063 => x"24fdea38",
  1064 => x"76802e94",
  1065 => x"3881ed52",
  1066 => x"b8f4519e",
  1067 => x"aa2db494",
  1068 => x"0852b8f4",
  1069 => x"519eaa2d",
  1070 => x"805372b2",
  1071 => x"e80c029c",
  1072 => x"050d0402",
  1073 => x"fc050d80",
  1074 => x"51800ba8",
  1075 => x"e81281b7",
  1076 => x"2d811151",
  1077 => x"81ff7125",
  1078 => x"f0380284",
  1079 => x"050d0402",
  1080 => x"f4050d74",
  1081 => x"51a29c2d",
  1082 => x"a8e81180",
  1083 => x"f52d7081",
  1084 => x"ff0671fd",
  1085 => x"06525452",
  1086 => x"71a8e812",
  1087 => x"81b72da2",
  1088 => x"962d72b2",
  1089 => x"e80c028c",
  1090 => x"050d0471",
  1091 => x"980c04ff",
  1092 => x"b008b2e8",
  1093 => x"0c04810b",
  1094 => x"ffb00c04",
  1095 => x"800bffb0",
  1096 => x"0c04b2f4",
  1097 => x"0802b2f4",
  1098 => x"0cff3d0d",
  1099 => x"800bb2f4",
  1100 => x"08fc050c",
  1101 => x"b2f40888",
  1102 => x"05088106",
  1103 => x"ff117009",
  1104 => x"70b2f408",
  1105 => x"8c050806",
  1106 => x"b2f408fc",
  1107 => x"050811b2",
  1108 => x"f408fc05",
  1109 => x"0cb2f408",
  1110 => x"88050881",
  1111 => x"2ab2f408",
  1112 => x"88050cb2",
  1113 => x"f4088c05",
  1114 => x"0810b2f4",
  1115 => x"088c050c",
  1116 => x"51515151",
  1117 => x"b2f40888",
  1118 => x"0508802e",
  1119 => x"8438ffb4",
  1120 => x"39b2f408",
  1121 => x"fc050870",
  1122 => x"b2e80c51",
  1123 => x"833d0db2",
  1124 => x"f40c0400",
  1125 => x"00ffffff",
  1126 => x"ff00ffff",
  1127 => x"ffff00ff",
  1128 => x"ffffff00",
  1129 => x"496e6974",
  1130 => x"69616c69",
  1131 => x"7a696e67",
  1132 => x"20534420",
  1133 => x"63617264",
  1134 => x"0a000000",
  1135 => x"48756e74",
  1136 => x"696e6720",
  1137 => x"666f7220",
  1138 => x"70617274",
  1139 => x"6974696f",
  1140 => x"6e0a0000",
  1141 => x"42494f53",
  1142 => x"5f4d3250",
  1143 => x"524f4d00",
  1144 => x"4f70656e",
  1145 => x"65642066",
  1146 => x"696c652c",
  1147 => x"206c6f61",
  1148 => x"64696e67",
  1149 => x"2e2e2e0a",
  1150 => x"00000000",
  1151 => x"52656164",
  1152 => x"20626c6f",
  1153 => x"636b2066",
  1154 => x"61696c65",
  1155 => x"640a0000",
  1156 => x"4c6f6164",
  1157 => x"696e6720",
  1158 => x"42494f53",
  1159 => x"20666169",
  1160 => x"6c65640a",
  1161 => x"00000000",
  1162 => x"496e6974",
  1163 => x"69616c69",
  1164 => x"73696e67",
  1165 => x"2050532f",
  1166 => x"3220696e",
  1167 => x"74657266",
  1168 => x"6163652e",
  1169 => x"2e2e0a00",
  1170 => x"52656164",
  1171 => x"696e6720",
  1172 => x"4d42520a",
  1173 => x"00000000",
  1174 => x"52656164",
  1175 => x"206f6620",
  1176 => x"4d425220",
  1177 => x"6661696c",
  1178 => x"65640a00",
  1179 => x"4d425220",
  1180 => x"73756363",
  1181 => x"65737366",
  1182 => x"756c6c79",
  1183 => x"20726561",
  1184 => x"640a0000",
  1185 => x"46415431",
  1186 => x"36202020",
  1187 => x"00000000",
  1188 => x"46415433",
  1189 => x"32202020",
  1190 => x"00000000",
  1191 => x"50617274",
  1192 => x"6974696f",
  1193 => x"6e636f75",
  1194 => x"6e742025",
  1195 => x"640a0000",
  1196 => x"4e6f2070",
  1197 => x"61727469",
  1198 => x"74696f6e",
  1199 => x"20736967",
  1200 => x"6e617475",
  1201 => x"72652066",
  1202 => x"6f756e64",
  1203 => x"0a000000",
  1204 => x"52656164",
  1205 => x"696e6720",
  1206 => x"626f6f74",
  1207 => x"20736563",
  1208 => x"746f7220",
  1209 => x"25640a00",
  1210 => x"52656164",
  1211 => x"20626f6f",
  1212 => x"74207365",
  1213 => x"63746f72",
  1214 => x"2066726f",
  1215 => x"6d206669",
  1216 => x"72737420",
  1217 => x"70617274",
  1218 => x"6974696f",
  1219 => x"6e0a0000",
  1220 => x"48756e74",
  1221 => x"696e6720",
  1222 => x"666f7220",
  1223 => x"66696c65",
  1224 => x"73797374",
  1225 => x"656d0a00",
  1226 => x"556e7375",
  1227 => x"70706f72",
  1228 => x"74656420",
  1229 => x"70617274",
  1230 => x"6974696f",
  1231 => x"6e207479",
  1232 => x"7065210d",
  1233 => x"00000000",
  1234 => x"436c7573",
  1235 => x"74657220",
  1236 => x"73697a65",
  1237 => x"3a202564",
  1238 => x"2c20436c",
  1239 => x"75737465",
  1240 => x"72206d61",
  1241 => x"736b2c20",
  1242 => x"25640a00",
  1243 => x"47657443",
  1244 => x"6c757374",
  1245 => x"65722072",
  1246 => x"65616469",
  1247 => x"6e672073",
  1248 => x"6563746f",
  1249 => x"72202564",
  1250 => x"0a000000",
  1251 => x"52656164",
  1252 => x"696e6720",
  1253 => x"64697265",
  1254 => x"63746f72",
  1255 => x"79207365",
  1256 => x"63746f72",
  1257 => x"2025640a",
  1258 => x"00000000",
  1259 => x"47657446",
  1260 => x"41544c69",
  1261 => x"6e6b2072",
  1262 => x"65747572",
  1263 => x"6e656420",
  1264 => x"25640a00",
  1265 => x"436d645f",
  1266 => x"696e6974",
  1267 => x"0a000000",
  1268 => x"636d645f",
  1269 => x"434d4438",
  1270 => x"20726573",
  1271 => x"706f6e73",
  1272 => x"653a2025",
  1273 => x"640a0000",
  1274 => x"434d4438",
  1275 => x"5f342072",
  1276 => x"6573706f",
  1277 => x"6e73653a",
  1278 => x"2025640a",
  1279 => x"00000000",
  1280 => x"53444843",
  1281 => x"20496e69",
  1282 => x"7469616c",
  1283 => x"697a6174",
  1284 => x"696f6e20",
  1285 => x"6572726f",
  1286 => x"72210a00",
  1287 => x"434d4435",
  1288 => x"38202564",
  1289 => x"0a202000",
  1290 => x"434d4435",
  1291 => x"385f3220",
  1292 => x"25640a20",
  1293 => x"20000000",
  1294 => x"53504920",
  1295 => x"496e6974",
  1296 => x"28290a00",
  1297 => x"52656164",
  1298 => x"20636f6d",
  1299 => x"6d616e64",
  1300 => x"20666169",
  1301 => x"6c656420",
  1302 => x"61742025",
  1303 => x"64202825",
  1304 => x"64290a00",
  1305 => x"ffffe000",
  1306 => x"00000000",
  1307 => x"00000000",
  1308 => x"00000000",
  1309 => x"00000000",
  1310 => x"00000000",
  1311 => x"00000000",
  1312 => x"00000000",
  1313 => x"00000000",
  1314 => x"00000000",
  1315 => x"00000000",
  1316 => x"00000000",
  1317 => x"00000000",
  1318 => x"00000000",
  1319 => x"00000000",
  1320 => x"00000000",
  1321 => x"00000000",
  1322 => x"00000000",
  1323 => x"00000000",
  1324 => x"00000000",
  1325 => x"00000000",
  1326 => x"00000000",
  1327 => x"00000000",
  1328 => x"00000000",
  1329 => x"00000000",
  1330 => x"00000000",
  1331 => x"00000000",
  1332 => x"00000000",
  1333 => x"00000000",
  1334 => x"00000000",
  1335 => x"00000000",
  1336 => x"00000000",
  1337 => x"00000000",
  1338 => x"00000000",
  1339 => x"00000000",
  1340 => x"00000000",
  1341 => x"00000000",
  1342 => x"00000000",
  1343 => x"00000000",
  1344 => x"00000000",
  1345 => x"00000000",
  1346 => x"00000000",
  1347 => x"00000000",
  1348 => x"00000000",
  1349 => x"00000000",
  1350 => x"00000000",
  1351 => x"00000000",
  1352 => x"00000000",
  1353 => x"00000000",
  1354 => x"00000000",
  1355 => x"00000000",
  1356 => x"00000000",
  1357 => x"00000000",
  1358 => x"00000000",
  1359 => x"00000000",
  1360 => x"00000000",
  1361 => x"00000000",
  1362 => x"00000000",
  1363 => x"00000000",
  1364 => x"00000000",
  1365 => x"00000000",
  1366 => x"00000000",
  1367 => x"00000000",
  1368 => x"00000000",
  1369 => x"00000000",
  1370 => x"00000000",
  1371 => x"00000000",
  1372 => x"00000000",
  1373 => x"00000000",
  1374 => x"00000000",
  1375 => x"00000000",
  1376 => x"00000000",
  1377 => x"00000000",
  1378 => x"00000000",
  1379 => x"00000000",
  1380 => x"00000000",
  1381 => x"00000000",
  1382 => x"00000000",
  1383 => x"00000009",
  1384 => x"00000000",
  1385 => x"00000000",
  1386 => x"00000000",
  1387 => x"00000000",
  1388 => x"00000000",
  1389 => x"00000000",
  1390 => x"00000000",
  1391 => x"00000071",
  1392 => x"00000031",
  1393 => x"00000000",
  1394 => x"00000000",
  1395 => x"00000000",
  1396 => x"0000007a",
  1397 => x"00000073",
  1398 => x"00000061",
  1399 => x"00000077",
  1400 => x"00000032",
  1401 => x"00000000",
  1402 => x"00000000",
  1403 => x"00000063",
  1404 => x"00000078",
  1405 => x"00000064",
  1406 => x"00000065",
  1407 => x"00000034",
  1408 => x"00000033",
  1409 => x"00000000",
  1410 => x"00000000",
  1411 => x"00000020",
  1412 => x"00000076",
  1413 => x"00000066",
  1414 => x"00000074",
  1415 => x"00000072",
  1416 => x"00000035",
  1417 => x"00000000",
  1418 => x"00000000",
  1419 => x"0000006e",
  1420 => x"00000062",
  1421 => x"00000068",
  1422 => x"00000067",
  1423 => x"00000079",
  1424 => x"00000036",
  1425 => x"00000000",
  1426 => x"00000000",
  1427 => x"00000000",
  1428 => x"0000006d",
  1429 => x"0000006a",
  1430 => x"00000075",
  1431 => x"00000037",
  1432 => x"00000038",
  1433 => x"00000000",
  1434 => x"00000000",
  1435 => x"0000002c",
  1436 => x"0000006b",
  1437 => x"00000069",
  1438 => x"0000006f",
  1439 => x"00000030",
  1440 => x"00000039",
  1441 => x"00000000",
  1442 => x"00000000",
  1443 => x"0000002e",
  1444 => x"0000002f",
  1445 => x"0000006c",
  1446 => x"0000003b",
  1447 => x"00000070",
  1448 => x"0000002d",
  1449 => x"00000000",
  1450 => x"00000000",
  1451 => x"00000000",
  1452 => x"00000027",
  1453 => x"00000000",
  1454 => x"0000005b",
  1455 => x"0000003d",
  1456 => x"00000000",
  1457 => x"00000000",
  1458 => x"00000000",
  1459 => x"00000000",
  1460 => x"0000000a",
  1461 => x"0000005d",
  1462 => x"00000000",
  1463 => x"00000023",
  1464 => x"00000000",
  1465 => x"00000000",
  1466 => x"00000000",
  1467 => x"00000000",
  1468 => x"00000000",
  1469 => x"00000000",
  1470 => x"00000000",
  1471 => x"00000000",
  1472 => x"00000008",
  1473 => x"00000000",
  1474 => x"00000000",
  1475 => x"00000031",
  1476 => x"00000000",
  1477 => x"00000034",
  1478 => x"00000037",
  1479 => x"00000000",
  1480 => x"00000000",
  1481 => x"00000000",
  1482 => x"00000030",
  1483 => x"0000002e",
  1484 => x"00000032",
  1485 => x"00000035",
  1486 => x"00000036",
  1487 => x"00000038",
  1488 => x"0000001b",
  1489 => x"00000000",
  1490 => x"00000000",
  1491 => x"0000002b",
  1492 => x"00000033",
  1493 => x"00000000",
  1494 => x"0000002a",
  1495 => x"00000039",
  1496 => x"00000000",
  1497 => x"00000000",
  1498 => x"00000000",
  1499 => x"00000000",
  1500 => x"00000000",
  1501 => x"00000000",
  1502 => x"00000000",
  1503 => x"00000000",
  1504 => x"00000000",
  1505 => x"00000000",
  1506 => x"00000000",
  1507 => x"00000000",
  1508 => x"00000000",
  1509 => x"00000000",
  1510 => x"00000000",
  1511 => x"00000008",
  1512 => x"00000000",
  1513 => x"00000000",
  1514 => x"00000000",
  1515 => x"00000000",
  1516 => x"00000000",
  1517 => x"00000000",
  1518 => x"00000000",
  1519 => x"00000051",
  1520 => x"00000021",
  1521 => x"00000000",
  1522 => x"00000000",
  1523 => x"00000000",
  1524 => x"0000005a",
  1525 => x"00000053",
  1526 => x"00000041",
  1527 => x"00000057",
  1528 => x"00000022",
  1529 => x"00000000",
  1530 => x"00000000",
  1531 => x"00000043",
  1532 => x"00000058",
  1533 => x"00000044",
  1534 => x"00000045",
  1535 => x"00000024",
  1536 => x"000000a3",
  1537 => x"00000000",
  1538 => x"00000000",
  1539 => x"00000020",
  1540 => x"00000056",
  1541 => x"00000046",
  1542 => x"00000054",
  1543 => x"00000052",
  1544 => x"00000025",
  1545 => x"00000000",
  1546 => x"00000000",
  1547 => x"0000004e",
  1548 => x"00000042",
  1549 => x"00000048",
  1550 => x"00000047",
  1551 => x"00000059",
  1552 => x"0000005e",
  1553 => x"00000000",
  1554 => x"00000000",
  1555 => x"00000000",
  1556 => x"0000004d",
  1557 => x"0000004a",
  1558 => x"00000055",
  1559 => x"00000026",
  1560 => x"0000002a",
  1561 => x"00000000",
  1562 => x"00000000",
  1563 => x"0000003c",
  1564 => x"0000004b",
  1565 => x"00000049",
  1566 => x"0000004f",
  1567 => x"00000029",
  1568 => x"00000028",
  1569 => x"00000000",
  1570 => x"00000000",
  1571 => x"0000003e",
  1572 => x"0000003f",
  1573 => x"0000004c",
  1574 => x"0000003a",
  1575 => x"00000050",
  1576 => x"0000005f",
  1577 => x"00000000",
  1578 => x"00000000",
  1579 => x"00000000",
  1580 => x"0000003f",
  1581 => x"00000000",
  1582 => x"0000007b",
  1583 => x"0000002b",
  1584 => x"00000000",
  1585 => x"00000000",
  1586 => x"00000000",
  1587 => x"00000000",
  1588 => x"0000000a",
  1589 => x"0000007d",
  1590 => x"00000000",
  1591 => x"0000007e",
  1592 => x"00000000",
  1593 => x"00000000",
  1594 => x"00000000",
  1595 => x"00000000",
  1596 => x"00000000",
  1597 => x"00000000",
  1598 => x"00000000",
  1599 => x"00000000",
  1600 => x"00000009",
  1601 => x"00000000",
  1602 => x"00000000",
  1603 => x"00000031",
  1604 => x"00000000",
  1605 => x"00000034",
  1606 => x"00000037",
  1607 => x"00000000",
  1608 => x"00000000",
  1609 => x"00000000",
  1610 => x"00000030",
  1611 => x"0000002e",
  1612 => x"00000032",
  1613 => x"00000035",
  1614 => x"00000036",
  1615 => x"00000038",
  1616 => x"0000001b",
  1617 => x"00000000",
  1618 => x"00000000",
  1619 => x"0000002b",
  1620 => x"00000033",
  1621 => x"00000000",
  1622 => x"0000002a",
  1623 => x"00000039",
  1624 => x"00000000",
  1625 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

