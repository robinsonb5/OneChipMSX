-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b0bb7",
     9 => x"ec080b0b",
    10 => x"0bb7f008",
    11 => x"0b0b0bb7",
    12 => x"f4080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"b7f40c0b",
    16 => x"0b0bb7f0",
    17 => x"0c0b0b0b",
    18 => x"b7ec0c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0baecc",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"b7ec70bd",
    57 => x"a4278b38",
    58 => x"80717084",
    59 => x"05530c81",
    60 => x"e2048c51",
    61 => x"8d8d0402",
    62 => x"fc050df8",
    63 => x"80518f0b",
    64 => x"b7fc0c9f",
    65 => x"0bb8800c",
    66 => x"a0717081",
    67 => x"055334b8",
    68 => x"8008ff05",
    69 => x"b8800cb8",
    70 => x"80088025",
    71 => x"eb38b7fc",
    72 => x"08ff05b7",
    73 => x"fc0cb7fc",
    74 => x"088025d7",
    75 => x"38028405",
    76 => x"0d0402f0",
    77 => x"050df880",
    78 => x"53f8a054",
    79 => x"83bf5273",
    80 => x"70810555",
    81 => x"33517073",
    82 => x"70810555",
    83 => x"34ff1252",
    84 => x"718025eb",
    85 => x"38fbc053",
    86 => x"9f52a073",
    87 => x"70810555",
    88 => x"34ff1252",
    89 => x"718025f2",
    90 => x"38029005",
    91 => x"0d0402f4",
    92 => x"050d7453",
    93 => x"8e0bb7fc",
    94 => x"08258f38",
    95 => x"82b22db7",
    96 => x"fc08ff05",
    97 => x"b7fc0c82",
    98 => x"f404b7fc",
    99 => x"08b88008",
   100 => x"5351728a",
   101 => x"2e098106",
   102 => x"b7387151",
   103 => x"719f24a0",
   104 => x"38b7fc08",
   105 => x"a02911f8",
   106 => x"80115151",
   107 => x"a07134b8",
   108 => x"80088105",
   109 => x"b8800cb8",
   110 => x"8008519f",
   111 => x"7125e238",
   112 => x"800bb880",
   113 => x"0cb7fc08",
   114 => x"8105b7fc",
   115 => x"0c83e404",
   116 => x"70a02912",
   117 => x"f8801151",
   118 => x"51727134",
   119 => x"b8800881",
   120 => x"05b8800c",
   121 => x"b88008a0",
   122 => x"2e098106",
   123 => x"8e38800b",
   124 => x"b8800cb7",
   125 => x"fc088105",
   126 => x"b7fc0c02",
   127 => x"8c050d04",
   128 => x"02e8050d",
   129 => x"77795656",
   130 => x"880bfc16",
   131 => x"77712c8f",
   132 => x"06545254",
   133 => x"80537272",
   134 => x"25953871",
   135 => x"53fbe014",
   136 => x"51877134",
   137 => x"8114ff14",
   138 => x"545472f1",
   139 => x"387153f9",
   140 => x"1576712c",
   141 => x"87065351",
   142 => x"71802e8b",
   143 => x"38fbe014",
   144 => x"51717134",
   145 => x"81145472",
   146 => x"8e249538",
   147 => x"8f733153",
   148 => x"fbe01451",
   149 => x"a0713481",
   150 => x"14ff1454",
   151 => x"5472f138",
   152 => x"0298050d",
   153 => x"0402ec05",
   154 => x"0d800bb8",
   155 => x"840cf68c",
   156 => x"08f69008",
   157 => x"71882c56",
   158 => x"5481ff06",
   159 => x"52737225",
   160 => x"88387154",
   161 => x"820bb884",
   162 => x"0c72882c",
   163 => x"7381ff06",
   164 => x"54557473",
   165 => x"258b3872",
   166 => x"b8840884",
   167 => x"07b8840c",
   168 => x"5573842b",
   169 => x"86a07125",
   170 => x"83713170",
   171 => x"0b0b0bb4",
   172 => x"cc0c8171",
   173 => x"2bff05f6",
   174 => x"880cfecc",
   175 => x"13ff122c",
   176 => x"788829ff",
   177 => x"94057081",
   178 => x"2cb88408",
   179 => x"52585255",
   180 => x"51525476",
   181 => x"802e8538",
   182 => x"70810751",
   183 => x"70f6940c",
   184 => x"71098105",
   185 => x"f6800c72",
   186 => x"098105f6",
   187 => x"840c0294",
   188 => x"050d0402",
   189 => x"f4050d74",
   190 => x"53727081",
   191 => x"055480f5",
   192 => x"2d527180",
   193 => x"2e893871",
   194 => x"5182ee2d",
   195 => x"85f90402",
   196 => x"8c050d04",
   197 => x"02f8050d",
   198 => x"a6822d80",
   199 => x"da51a7b9",
   200 => x"2db7ec08",
   201 => x"812a7081",
   202 => x"06515271",
   203 => x"802ee938",
   204 => x"0288050d",
   205 => x"0402f405",
   206 => x"0dbd9408",
   207 => x"99c406b6",
   208 => x"c80b80f5",
   209 => x"2d525270",
   210 => x"802e8638",
   211 => x"71848007",
   212 => x"52b6800b",
   213 => x"80f52d72",
   214 => x"07b6a40b",
   215 => x"80f52d70",
   216 => x"812a7081",
   217 => x"06515354",
   218 => x"5270802e",
   219 => x"86387182",
   220 => x"80075272",
   221 => x"81065170",
   222 => x"802e8538",
   223 => x"71880752",
   224 => x"b6b00b80",
   225 => x"f52d7084",
   226 => x"2b730781",
   227 => x"8432b7ec",
   228 => x"0c51028c",
   229 => x"050d0402",
   230 => x"f4050d74",
   231 => x"70818432",
   232 => x"bd940c70",
   233 => x"83065253",
   234 => x"70b5f80b",
   235 => x"880581b7",
   236 => x"2d72892a",
   237 => x"70810651",
   238 => x"5170b6c8",
   239 => x"0b81b72d",
   240 => x"72832a81",
   241 => x"0673882a",
   242 => x"70810651",
   243 => x"52527080",
   244 => x"2e853871",
   245 => x"82075271",
   246 => x"b6a40b81",
   247 => x"b72d7284",
   248 => x"2c708306",
   249 => x"515170b6",
   250 => x"b00b81b7",
   251 => x"2d70b7ec",
   252 => x"0c028c05",
   253 => x"0d0402f4",
   254 => x"050db5b0",
   255 => x"0b881180",
   256 => x"f52d8c12",
   257 => x"881180f5",
   258 => x"2d70842b",
   259 => x"73078c13",
   260 => x"881180f5",
   261 => x"2d70882b",
   262 => x"73079413",
   263 => x"80f52d70",
   264 => x"8c2b7207",
   265 => x"b7ec0c53",
   266 => x"53535353",
   267 => x"56525351",
   268 => x"028c050d",
   269 => x"0402f405",
   270 => x"0d74b5b0",
   271 => x"71870655",
   272 => x"53517288",
   273 => x"1381b72d",
   274 => x"8c127184",
   275 => x"2c708706",
   276 => x"55525272",
   277 => x"881381b7",
   278 => x"2d8c1271",
   279 => x"842c7087",
   280 => x"06555252",
   281 => x"72881381",
   282 => x"b72d7084",
   283 => x"2c708706",
   284 => x"51517094",
   285 => x"1381b72d",
   286 => x"028c050d",
   287 => x"0402d405",
   288 => x"0db1cc51",
   289 => x"85f32d9d",
   290 => x"b32db7ec",
   291 => x"08802e83",
   292 => x"a23886b5",
   293 => x"2db7ec08",
   294 => x"538ffc2d",
   295 => x"b7ec0854",
   296 => x"b7ec0880",
   297 => x"2e838e38",
   298 => x"a1b62db7",
   299 => x"ec08802e",
   300 => x"8738b1e4",
   301 => x"5189c504",
   302 => x"999f2db7",
   303 => x"ec08802e",
   304 => x"a238b1f8",
   305 => x"5185f32d",
   306 => x"b2905185",
   307 => x"f32d8694",
   308 => x"2d728407",
   309 => x"53810bfe",
   310 => x"c40c72fe",
   311 => x"c00c7251",
   312 => x"87972d84",
   313 => x"0bfec40c",
   314 => x"b2ac52b8",
   315 => x"8c51968e",
   316 => x"2db7ec08",
   317 => x"802e80e1",
   318 => x"387c802e",
   319 => x"af3872b8",
   320 => x"980c87f6",
   321 => x"2db7ec08",
   322 => x"b89c0cb8",
   323 => x"a05480fd",
   324 => x"53807470",
   325 => x"8405560c",
   326 => x"ff135372",
   327 => x"8025f238",
   328 => x"b89852b8",
   329 => x"8c5198f9",
   330 => x"2d8ad904",
   331 => x"b2ac52b8",
   332 => x"8c51968e",
   333 => x"2db7ec08",
   334 => x"802e9e38",
   335 => x"b89852b8",
   336 => x"8c5198d3",
   337 => x"2db89808",
   338 => x"b89c0852",
   339 => x"5388b52d",
   340 => x"72fec00c",
   341 => x"72518797",
   342 => x"2db2b851",
   343 => x"85f32db2",
   344 => x"d052b88c",
   345 => x"51968e2d",
   346 => x"b7ec0898",
   347 => x"38b2dc51",
   348 => x"85f32db2",
   349 => x"f452b88c",
   350 => x"51968e2d",
   351 => x"b7ec0880",
   352 => x"2e81b038",
   353 => x"b3805185",
   354 => x"f32db890",
   355 => x"08578077",
   356 => x"595a767a",
   357 => x"2e8b3881",
   358 => x"1a78812a",
   359 => x"595a77f7",
   360 => x"38f71a5a",
   361 => x"80772581",
   362 => x"80387952",
   363 => x"77518480",
   364 => x"2db89852",
   365 => x"b88c5198",
   366 => x"d32db7ec",
   367 => x"0853b7ec",
   368 => x"08802e80",
   369 => x"c938b898",
   370 => x"5b80598b",
   371 => x"fb047a70",
   372 => x"84055c08",
   373 => x"7081ff06",
   374 => x"71882c70",
   375 => x"81ff0673",
   376 => x"902c7081",
   377 => x"ff067598",
   378 => x"2afec80c",
   379 => x"fec80c58",
   380 => x"fec80c57",
   381 => x"fec80c84",
   382 => x"1a5a5376",
   383 => x"53848077",
   384 => x"25843884",
   385 => x"80537279",
   386 => x"24c4388c",
   387 => x"9904b390",
   388 => x"5185f32d",
   389 => x"72548cb5",
   390 => x"04b88c51",
   391 => x"98a62dfc",
   392 => x"80178119",
   393 => x"59578ba4",
   394 => x"04820bfe",
   395 => x"c40c8154",
   396 => x"8cb50480",
   397 => x"5473b7ec",
   398 => x"0c02ac05",
   399 => x"0d0402f8",
   400 => x"050da889",
   401 => x"2d81f72d",
   402 => x"815184e5",
   403 => x"2dfec452",
   404 => x"81720ca5",
   405 => x"822da582",
   406 => x"2d84720c",
   407 => x"735188fd",
   408 => x"2db4d051",
   409 => x"a9e72d80",
   410 => x"5184e52d",
   411 => x"0288050d",
   412 => x"0402fc05",
   413 => x"0d81518c",
   414 => x"be2d0284",
   415 => x"050d0402",
   416 => x"fc050d80",
   417 => x"518cbe2d",
   418 => x"0284050d",
   419 => x"0402ec05",
   420 => x"0d84b851",
   421 => x"87972d81",
   422 => x"0bfec40c",
   423 => x"84b80bfe",
   424 => x"c00c840b",
   425 => x"fec40c83",
   426 => x"0bfecc0c",
   427 => x"a59d2da7",
   428 => x"fd2da582",
   429 => x"2da5822d",
   430 => x"81f72d81",
   431 => x"5184e52d",
   432 => x"a5822da5",
   433 => x"822d8151",
   434 => x"84e52d80",
   435 => x"5188fd2d",
   436 => x"b7ec0880",
   437 => x"2e81d238",
   438 => x"805184e5",
   439 => x"2db4d051",
   440 => x"a9e72dbc",
   441 => x"f4088938",
   442 => x"bcf80880",
   443 => x"2e80e238",
   444 => x"fed00870",
   445 => x"81065152",
   446 => x"71802e80",
   447 => x"d438a883",
   448 => x"2dbcf408",
   449 => x"70bcf808",
   450 => x"70575556",
   451 => x"5280ff72",
   452 => x"25843880",
   453 => x"ff5280ff",
   454 => x"73258438",
   455 => x"80ff5371",
   456 => x"ff802584",
   457 => x"38ff8052",
   458 => x"72ff8025",
   459 => x"8438ff80",
   460 => x"53747231",
   461 => x"bcf40c73",
   462 => x"7331bcf8",
   463 => x"0ca7fd2d",
   464 => x"71882b83",
   465 => x"fe800673",
   466 => x"81ff0671",
   467 => x"07fed00c",
   468 => x"52a6822d",
   469 => x"a9f72db7",
   470 => x"ec085386",
   471 => x"b52db7ec",
   472 => x"08fec00c",
   473 => x"87f62db7",
   474 => x"ec08fed4",
   475 => x"0c86b52d",
   476 => x"b7ec08b8",
   477 => x"88082e9c",
   478 => x"38b7ec08",
   479 => x"b8880c84",
   480 => x"52725184",
   481 => x"e52da582",
   482 => x"2da5822d",
   483 => x"ff125271",
   484 => x"8025ee38",
   485 => x"72802e89",
   486 => x"388a0bfe",
   487 => x"c40c8de3",
   488 => x"04820bfe",
   489 => x"c40c8de3",
   490 => x"04b3a051",
   491 => x"85f32d82",
   492 => x"0bfec40c",
   493 => x"800bb7ec",
   494 => x"0c029405",
   495 => x"0d0402e8",
   496 => x"050d7779",
   497 => x"7b585555",
   498 => x"80537276",
   499 => x"25a33874",
   500 => x"70810556",
   501 => x"80f52d74",
   502 => x"70810556",
   503 => x"80f52d52",
   504 => x"5271712e",
   505 => x"86388151",
   506 => x"8ff30481",
   507 => x"13538fca",
   508 => x"04805170",
   509 => x"b7ec0c02",
   510 => x"98050d04",
   511 => x"02d8050d",
   512 => x"800bbca0",
   513 => x"0cb89852",
   514 => x"8051a09b",
   515 => x"2db7ec08",
   516 => x"54b7ec08",
   517 => x"8c38b3b8",
   518 => x"5185f32d",
   519 => x"73559597",
   520 => x"04805681",
   521 => x"0bbcc40c",
   522 => x"8853b3c4",
   523 => x"52b8ce51",
   524 => x"8fbe2db7",
   525 => x"ec08762e",
   526 => x"09810687",
   527 => x"38b7ec08",
   528 => x"bcc40c88",
   529 => x"53b3d052",
   530 => x"b8ea518f",
   531 => x"be2db7ec",
   532 => x"088738b7",
   533 => x"ec08bcc4",
   534 => x"0cbcc408",
   535 => x"802e80f6",
   536 => x"38bbde0b",
   537 => x"80f52dbb",
   538 => x"df0b80f5",
   539 => x"2d71982b",
   540 => x"71902b07",
   541 => x"bbe00b80",
   542 => x"f52d7088",
   543 => x"2b7207bb",
   544 => x"e10b80f5",
   545 => x"2d7107bc",
   546 => x"960b80f5",
   547 => x"2dbc970b",
   548 => x"80f52d71",
   549 => x"882b0753",
   550 => x"5f54525a",
   551 => x"56575573",
   552 => x"81abaa2e",
   553 => x"0981068d",
   554 => x"387551a1",
   555 => x"bd2db7ec",
   556 => x"085691c2",
   557 => x"047382d4",
   558 => x"d52e8738",
   559 => x"b3dc5192",
   560 => x"8304b898",
   561 => x"527551a0",
   562 => x"9b2db7ec",
   563 => x"0855b7ec",
   564 => x"08802e83",
   565 => x"c2388853",
   566 => x"b3d052b8",
   567 => x"ea518fbe",
   568 => x"2db7ec08",
   569 => x"8938810b",
   570 => x"bca00c92",
   571 => x"89048853",
   572 => x"b3c452b8",
   573 => x"ce518fbe",
   574 => x"2db7ec08",
   575 => x"802e8a38",
   576 => x"b3f05185",
   577 => x"f32d92e3",
   578 => x"04bc960b",
   579 => x"80f52d54",
   580 => x"7380d52e",
   581 => x"09810680",
   582 => x"ca38bc97",
   583 => x"0b80f52d",
   584 => x"547381aa",
   585 => x"2e098106",
   586 => x"ba38800b",
   587 => x"b8980b80",
   588 => x"f52d5654",
   589 => x"7481e92e",
   590 => x"83388154",
   591 => x"7481eb2e",
   592 => x"8c388055",
   593 => x"73752e09",
   594 => x"810682cb",
   595 => x"38b8a30b",
   596 => x"80f52d55",
   597 => x"748d38b8",
   598 => x"a40b80f5",
   599 => x"2d547382",
   600 => x"2e863880",
   601 => x"55959704",
   602 => x"b8a50b80",
   603 => x"f52d70bc",
   604 => x"980cff05",
   605 => x"bc9c0cb8",
   606 => x"a60b80f5",
   607 => x"2db8a70b",
   608 => x"80f52d58",
   609 => x"76057782",
   610 => x"80290570",
   611 => x"bca40cb8",
   612 => x"a80b80f5",
   613 => x"2d70bcb8",
   614 => x"0cbca008",
   615 => x"59575876",
   616 => x"802e81a3",
   617 => x"388853b3",
   618 => x"d052b8ea",
   619 => x"518fbe2d",
   620 => x"b7ec0881",
   621 => x"e238bc98",
   622 => x"0870842b",
   623 => x"bcbc0c70",
   624 => x"bcb40cb8",
   625 => x"bd0b80f5",
   626 => x"2db8bc0b",
   627 => x"80f52d71",
   628 => x"82802905",
   629 => x"b8be0b80",
   630 => x"f52d7084",
   631 => x"80802912",
   632 => x"b8bf0b80",
   633 => x"f52d7081",
   634 => x"800a2912",
   635 => x"70bcc00c",
   636 => x"bcb80871",
   637 => x"29bca408",
   638 => x"0570bca8",
   639 => x"0cb8c50b",
   640 => x"80f52db8",
   641 => x"c40b80f5",
   642 => x"2d718280",
   643 => x"2905b8c6",
   644 => x"0b80f52d",
   645 => x"70848080",
   646 => x"2912b8c7",
   647 => x"0b80f52d",
   648 => x"70982b81",
   649 => x"f00a0672",
   650 => x"0570bcac",
   651 => x"0cfe117e",
   652 => x"297705bc",
   653 => x"b00c5259",
   654 => x"5243545e",
   655 => x"51525952",
   656 => x"5d575957",
   657 => x"959504b8",
   658 => x"aa0b80f5",
   659 => x"2db8a90b",
   660 => x"80f52d71",
   661 => x"82802905",
   662 => x"70bcbc0c",
   663 => x"70a02983",
   664 => x"ff057089",
   665 => x"2a70bcb4",
   666 => x"0cb8af0b",
   667 => x"80f52db8",
   668 => x"ae0b80f5",
   669 => x"2d718280",
   670 => x"290570bc",
   671 => x"c00c7b71",
   672 => x"291e70bc",
   673 => x"b00c7dbc",
   674 => x"ac0c7305",
   675 => x"bca80c55",
   676 => x"5e515155",
   677 => x"55815574",
   678 => x"b7ec0c02",
   679 => x"a8050d04",
   680 => x"02ec050d",
   681 => x"7670872c",
   682 => x"7180ff06",
   683 => x"555654bc",
   684 => x"a0088a38",
   685 => x"73882c74",
   686 => x"81ff0654",
   687 => x"55b89852",
   688 => x"bca40815",
   689 => x"51a09b2d",
   690 => x"b7ec0854",
   691 => x"b7ec0880",
   692 => x"2eb338bc",
   693 => x"a008802e",
   694 => x"98387284",
   695 => x"29b89805",
   696 => x"70085253",
   697 => x"a1bd2db7",
   698 => x"ec08f00a",
   699 => x"06539683",
   700 => x"047210b8",
   701 => x"98057080",
   702 => x"e02d5253",
   703 => x"a1ed2db7",
   704 => x"ec085372",
   705 => x"5473b7ec",
   706 => x"0c029405",
   707 => x"0d0402c8",
   708 => x"050d7f61",
   709 => x"5f5b800b",
   710 => x"bcac08bc",
   711 => x"b008595d",
   712 => x"56bca008",
   713 => x"762e8a38",
   714 => x"bc980884",
   715 => x"2b5896b7",
   716 => x"04bcb408",
   717 => x"842b5880",
   718 => x"59787827",
   719 => x"81a93878",
   720 => x"8f06a017",
   721 => x"5754738f",
   722 => x"38b89852",
   723 => x"76518117",
   724 => x"57a09b2d",
   725 => x"b8985680",
   726 => x"7680f52d",
   727 => x"56547474",
   728 => x"2e833881",
   729 => x"547481e5",
   730 => x"2e80f638",
   731 => x"81707506",
   732 => x"555d7380",
   733 => x"2e80ea38",
   734 => x"8b1680f5",
   735 => x"2d98065a",
   736 => x"7980de38",
   737 => x"8b537d52",
   738 => x"75518fbe",
   739 => x"2db7ec08",
   740 => x"80cf389c",
   741 => x"160851a1",
   742 => x"bd2db7ec",
   743 => x"08841c0c",
   744 => x"9a1680e0",
   745 => x"2d51a1ed",
   746 => x"2db7ec08",
   747 => x"b7ec0888",
   748 => x"1d0cb7ec",
   749 => x"085555bc",
   750 => x"a008802e",
   751 => x"98389416",
   752 => x"80e02d51",
   753 => x"a1ed2db7",
   754 => x"ec08902b",
   755 => x"83fff00a",
   756 => x"06701651",
   757 => x"5473881c",
   758 => x"0c797b0c",
   759 => x"7c54989d",
   760 => x"04811959",
   761 => x"96b904bc",
   762 => x"a008802e",
   763 => x"ae387b51",
   764 => x"95a02db7",
   765 => x"ec08b7ec",
   766 => x"0880ffff",
   767 => x"fff80655",
   768 => x"5c7380ff",
   769 => x"fffff82e",
   770 => x"9238b7ec",
   771 => x"08fe05bc",
   772 => x"980829bc",
   773 => x"a8080557",
   774 => x"96b70480",
   775 => x"5473b7ec",
   776 => x"0c02b805",
   777 => x"0d0402f4",
   778 => x"050d7470",
   779 => x"08810571",
   780 => x"0c7008bc",
   781 => x"9c080653",
   782 => x"53718e38",
   783 => x"88130851",
   784 => x"95a02db7",
   785 => x"ec088814",
   786 => x"0c810bb7",
   787 => x"ec0c028c",
   788 => x"050d0402",
   789 => x"f0050d75",
   790 => x"881108fe",
   791 => x"05bc9808",
   792 => x"29bca808",
   793 => x"117208bc",
   794 => x"9c080605",
   795 => x"79555354",
   796 => x"54a09b2d",
   797 => x"0290050d",
   798 => x"0402f005",
   799 => x"0d758811",
   800 => x"08fe05bc",
   801 => x"980829bc",
   802 => x"a8081172",
   803 => x"08bc9c08",
   804 => x"06057955",
   805 => x"5354549e",
   806 => x"db2d0290",
   807 => x"050d04bc",
   808 => x"a008b7ec",
   809 => x"0c0402f4",
   810 => x"050dd452",
   811 => x"81ff720c",
   812 => x"71085381",
   813 => x"ff720c72",
   814 => x"882b83fe",
   815 => x"80067208",
   816 => x"7081ff06",
   817 => x"51525381",
   818 => x"ff720c72",
   819 => x"7107882b",
   820 => x"72087081",
   821 => x"ff065152",
   822 => x"5381ff72",
   823 => x"0c727107",
   824 => x"882b7208",
   825 => x"7081ff06",
   826 => x"7207b7ec",
   827 => x"0c525302",
   828 => x"8c050d04",
   829 => x"02f4050d",
   830 => x"74767181",
   831 => x"ff06d40c",
   832 => x"5353bcc8",
   833 => x"08853871",
   834 => x"892b5271",
   835 => x"982ad40c",
   836 => x"71902a70",
   837 => x"81ff06d4",
   838 => x"0c517188",
   839 => x"2a7081ff",
   840 => x"06d40c51",
   841 => x"7181ff06",
   842 => x"d40c7290",
   843 => x"2a7081ff",
   844 => x"06d40c51",
   845 => x"d4087081",
   846 => x"ff065151",
   847 => x"82b8bf52",
   848 => x"7081ff2e",
   849 => x"09810694",
   850 => x"3881ff0b",
   851 => x"d40cd408",
   852 => x"7081ff06",
   853 => x"ff145451",
   854 => x"5171e538",
   855 => x"70b7ec0c",
   856 => x"028c050d",
   857 => x"0402fc05",
   858 => x"0d81c751",
   859 => x"81ff0bd4",
   860 => x"0cff1151",
   861 => x"708025f4",
   862 => x"38028405",
   863 => x"0d0402f0",
   864 => x"050d9ae5",
   865 => x"2d8fcf53",
   866 => x"805287fc",
   867 => x"80f75199",
   868 => x"f42db7ec",
   869 => x"0854b7ec",
   870 => x"08812e09",
   871 => x"8106a338",
   872 => x"81ff0bd4",
   873 => x"0c820a52",
   874 => x"849c80e9",
   875 => x"5199f42d",
   876 => x"b7ec088b",
   877 => x"3881ff0b",
   878 => x"d40c7353",
   879 => x"9bc8049a",
   880 => x"e52dff13",
   881 => x"5372c138",
   882 => x"72b7ec0c",
   883 => x"0290050d",
   884 => x"0402f405",
   885 => x"0d81ff0b",
   886 => x"d40c9353",
   887 => x"805287fc",
   888 => x"80c15199",
   889 => x"f42db7ec",
   890 => x"088b3881",
   891 => x"ff0bd40c",
   892 => x"81539bfe",
   893 => x"049ae52d",
   894 => x"ff135372",
   895 => x"df3872b7",
   896 => x"ec0c028c",
   897 => x"050d0402",
   898 => x"f0050d9a",
   899 => x"e52d83aa",
   900 => x"52849c80",
   901 => x"c85199f4",
   902 => x"2db7ec08",
   903 => x"812e0981",
   904 => x"06923899",
   905 => x"a62db7ec",
   906 => x"0883ffff",
   907 => x"06537283",
   908 => x"aa2e9738",
   909 => x"9bd12d9c",
   910 => x"c5048154",
   911 => x"9daa04b3",
   912 => x"fc5185f3",
   913 => x"2d80549d",
   914 => x"aa0481ff",
   915 => x"0bd40cb1",
   916 => x"539afe2d",
   917 => x"b7ec0880",
   918 => x"2e80c038",
   919 => x"805287fc",
   920 => x"80fa5199",
   921 => x"f42db7ec",
   922 => x"08b13881",
   923 => x"ff0bd40c",
   924 => x"d4085381",
   925 => x"ff0bd40c",
   926 => x"81ff0bd4",
   927 => x"0c81ff0b",
   928 => x"d40c81ff",
   929 => x"0bd40c72",
   930 => x"862a7081",
   931 => x"06b7ec08",
   932 => x"56515372",
   933 => x"802e9338",
   934 => x"9cba0472",
   935 => x"822eff9f",
   936 => x"38ff1353",
   937 => x"72ffaa38",
   938 => x"725473b7",
   939 => x"ec0c0290",
   940 => x"050d0402",
   941 => x"f0050d81",
   942 => x"0bbcc80c",
   943 => x"8454d008",
   944 => x"708f2a70",
   945 => x"81065151",
   946 => x"5372f338",
   947 => x"72d00c9a",
   948 => x"e52db48c",
   949 => x"5185f32d",
   950 => x"d008708f",
   951 => x"2a708106",
   952 => x"51515372",
   953 => x"f338810b",
   954 => x"d00cb153",
   955 => x"805284d4",
   956 => x"80c05199",
   957 => x"f42db7ec",
   958 => x"08812ea1",
   959 => x"3872822e",
   960 => x"0981068c",
   961 => x"38b49851",
   962 => x"85f32d80",
   963 => x"539ed204",
   964 => x"ff135372",
   965 => x"d738ff14",
   966 => x"5473ffa2",
   967 => x"389c872d",
   968 => x"b7ec08bc",
   969 => x"c80cb7ec",
   970 => x"088b3881",
   971 => x"5287fc80",
   972 => x"d05199f4",
   973 => x"2d81ff0b",
   974 => x"d40cd008",
   975 => x"708f2a70",
   976 => x"81065151",
   977 => x"5372f338",
   978 => x"72d00c81",
   979 => x"ff0bd40c",
   980 => x"815372b7",
   981 => x"ec0c0290",
   982 => x"050d0402",
   983 => x"e8050d78",
   984 => x"5681ff0b",
   985 => x"d40cd008",
   986 => x"708f2a70",
   987 => x"81065151",
   988 => x"5372f338",
   989 => x"82810bd0",
   990 => x"0c81ff0b",
   991 => x"d40c7752",
   992 => x"87fc80d8",
   993 => x"5199f42d",
   994 => x"b7ec0880",
   995 => x"2e8c38b4",
   996 => x"b05185f3",
   997 => x"2d8153a0",
   998 => x"920481ff",
   999 => x"0bd40c81",
  1000 => x"fe0bd40c",
  1001 => x"80ff5575",
  1002 => x"70840557",
  1003 => x"0870982a",
  1004 => x"d40c7090",
  1005 => x"2c7081ff",
  1006 => x"06d40c54",
  1007 => x"70882c70",
  1008 => x"81ff06d4",
  1009 => x"0c547081",
  1010 => x"ff06d40c",
  1011 => x"54ff1555",
  1012 => x"748025d3",
  1013 => x"3881ff0b",
  1014 => x"d40c81ff",
  1015 => x"0bd40c81",
  1016 => x"ff0bd40c",
  1017 => x"868da054",
  1018 => x"81ff0bd4",
  1019 => x"0cd40881",
  1020 => x"ff065574",
  1021 => x"8738ff14",
  1022 => x"5473ed38",
  1023 => x"81ff0bd4",
  1024 => x"0cd00870",
  1025 => x"8f2a7081",
  1026 => x"06515153",
  1027 => x"72f33872",
  1028 => x"d00c72b7",
  1029 => x"ec0c0298",
  1030 => x"050d0402",
  1031 => x"e8050d78",
  1032 => x"55805681",
  1033 => x"ff0bd40c",
  1034 => x"d008708f",
  1035 => x"2a708106",
  1036 => x"51515372",
  1037 => x"f3388281",
  1038 => x"0bd00c81",
  1039 => x"ff0bd40c",
  1040 => x"775287fc",
  1041 => x"80d15199",
  1042 => x"f42d80db",
  1043 => x"c6df54b7",
  1044 => x"ec08802e",
  1045 => x"8a38b390",
  1046 => x"5185f32d",
  1047 => x"a1ad0481",
  1048 => x"ff0bd40c",
  1049 => x"d4087081",
  1050 => x"ff065153",
  1051 => x"7281fe2e",
  1052 => x"0981069d",
  1053 => x"3880ff53",
  1054 => x"99a62db7",
  1055 => x"ec087570",
  1056 => x"8405570c",
  1057 => x"ff135372",
  1058 => x"8025ed38",
  1059 => x"8156a197",
  1060 => x"04ff1454",
  1061 => x"73c93881",
  1062 => x"ff0bd40c",
  1063 => x"d008708f",
  1064 => x"2a708106",
  1065 => x"51515372",
  1066 => x"f33872d0",
  1067 => x"0c75b7ec",
  1068 => x"0c029805",
  1069 => x"0d04bcc8",
  1070 => x"08b7ec0c",
  1071 => x"0402f405",
  1072 => x"0d747088",
  1073 => x"2a83fe80",
  1074 => x"06707298",
  1075 => x"2a077288",
  1076 => x"2b87fc80",
  1077 => x"80067398",
  1078 => x"2b81f00a",
  1079 => x"06717307",
  1080 => x"07b7ec0c",
  1081 => x"56515351",
  1082 => x"028c050d",
  1083 => x"0402f805",
  1084 => x"0d028e05",
  1085 => x"80f52d74",
  1086 => x"882b0770",
  1087 => x"83ffff06",
  1088 => x"b7ec0c51",
  1089 => x"0288050d",
  1090 => x"0402fc05",
  1091 => x"0d725180",
  1092 => x"710c800b",
  1093 => x"84120c02",
  1094 => x"84050d04",
  1095 => x"02f0050d",
  1096 => x"75700884",
  1097 => x"12085353",
  1098 => x"53ff5471",
  1099 => x"712ea838",
  1100 => x"a8832d84",
  1101 => x"13087084",
  1102 => x"29148811",
  1103 => x"70087081",
  1104 => x"ff068418",
  1105 => x"08811187",
  1106 => x"06841a0c",
  1107 => x"53515551",
  1108 => x"5151a7fd",
  1109 => x"2d715473",
  1110 => x"b7ec0c02",
  1111 => x"90050d04",
  1112 => x"02f4050d",
  1113 => x"a8832de0",
  1114 => x"08e40871",
  1115 => x"8b2a7081",
  1116 => x"06515354",
  1117 => x"5270802e",
  1118 => x"9d38bccc",
  1119 => x"08708429",
  1120 => x"bcd40573",
  1121 => x"81ff0671",
  1122 => x"0c5151bc",
  1123 => x"cc088111",
  1124 => x"8706bccc",
  1125 => x"0c51728b",
  1126 => x"2a708106",
  1127 => x"51517080",
  1128 => x"2e819238",
  1129 => x"b79c0884",
  1130 => x"29bd8005",
  1131 => x"7381ff06",
  1132 => x"710c51b7",
  1133 => x"9c088105",
  1134 => x"b79c0c85",
  1135 => x"0bb7980c",
  1136 => x"b79c08b7",
  1137 => x"94082e09",
  1138 => x"810681a6",
  1139 => x"38800bb7",
  1140 => x"9c0cbd90",
  1141 => x"08819b38",
  1142 => x"bd800870",
  1143 => x"09708306",
  1144 => x"fecc0c52",
  1145 => x"70852a70",
  1146 => x"8106bcf8",
  1147 => x"08555152",
  1148 => x"5370802e",
  1149 => x"8e38bd88",
  1150 => x"08fe8032",
  1151 => x"12bcf80c",
  1152 => x"a48a04bd",
  1153 => x"880812bc",
  1154 => x"f80c7284",
  1155 => x"2a708106",
  1156 => x"bcf40854",
  1157 => x"51517080",
  1158 => x"2e9038bd",
  1159 => x"840881ff",
  1160 => x"32128105",
  1161 => x"bcf40ca4",
  1162 => x"f20471bd",
  1163 => x"840831bc",
  1164 => x"f40ca4f2",
  1165 => x"04b79808",
  1166 => x"ff05b798",
  1167 => x"0cb79808",
  1168 => x"ff2e0981",
  1169 => x"06ac38b7",
  1170 => x"9c08802e",
  1171 => x"9238810b",
  1172 => x"bd900c87",
  1173 => x"0bb79408",
  1174 => x"31b7940c",
  1175 => x"a4ed04bd",
  1176 => x"90085170",
  1177 => x"802e8638",
  1178 => x"ff11bd90",
  1179 => x"0c800bb7",
  1180 => x"9c0c800b",
  1181 => x"bcfc0ca7",
  1182 => x"f62da7fd",
  1183 => x"2d028c05",
  1184 => x"0d0402fc",
  1185 => x"050da883",
  1186 => x"2d810bbc",
  1187 => x"fc0ca7fd",
  1188 => x"2dbcfc08",
  1189 => x"5170fa38",
  1190 => x"0284050d",
  1191 => x"0402f805",
  1192 => x"0dbccc51",
  1193 => x"a2892d80",
  1194 => x"0bbd900c",
  1195 => x"830bb794",
  1196 => x"0ce40870",
  1197 => x"8c2a7081",
  1198 => x"06515152",
  1199 => x"71802e86",
  1200 => x"38840bb7",
  1201 => x"940ce408",
  1202 => x"708d2a70",
  1203 => x"81065151",
  1204 => x"5271802e",
  1205 => x"9f38870b",
  1206 => x"b7940831",
  1207 => x"b7940ce4",
  1208 => x"08708a2a",
  1209 => x"70810651",
  1210 => x"51527180",
  1211 => x"2ef13881",
  1212 => x"f40be40c",
  1213 => x"a2e051a7",
  1214 => x"f22da79c",
  1215 => x"2d028805",
  1216 => x"0d0402f4",
  1217 => x"050da784",
  1218 => x"04b7ec08",
  1219 => x"81f02e09",
  1220 => x"81068938",
  1221 => x"810bb7e0",
  1222 => x"0ca78404",
  1223 => x"b7ec0881",
  1224 => x"e02e0981",
  1225 => x"06893881",
  1226 => x"0bb7e40c",
  1227 => x"a78404b7",
  1228 => x"ec0852b7",
  1229 => x"e408802e",
  1230 => x"8838b7ec",
  1231 => x"08818005",
  1232 => x"5271842c",
  1233 => x"728f0653",
  1234 => x"53b7e008",
  1235 => x"802e9938",
  1236 => x"728429b7",
  1237 => x"a0057213",
  1238 => x"81712b70",
  1239 => x"09730806",
  1240 => x"730c5153",
  1241 => x"53a6fa04",
  1242 => x"728429b7",
  1243 => x"a0057213",
  1244 => x"83712b72",
  1245 => x"0807720c",
  1246 => x"5353800b",
  1247 => x"b7e40c80",
  1248 => x"0bb7e00c",
  1249 => x"bccc51a2",
  1250 => x"9c2db7ec",
  1251 => x"08ff24fe",
  1252 => x"f838800b",
  1253 => x"b7ec0c02",
  1254 => x"8c050d04",
  1255 => x"02f8050d",
  1256 => x"b7a0528f",
  1257 => x"51807270",
  1258 => x"8405540c",
  1259 => x"ff115170",
  1260 => x"8025f238",
  1261 => x"0288050d",
  1262 => x"0402f005",
  1263 => x"0d7551a8",
  1264 => x"832d7082",
  1265 => x"2cfc06b7",
  1266 => x"a0117210",
  1267 => x"9e067108",
  1268 => x"70722a70",
  1269 => x"83068274",
  1270 => x"2b700974",
  1271 => x"06760c54",
  1272 => x"51565753",
  1273 => x"5153a7fd",
  1274 => x"2d71b7ec",
  1275 => x"0c029005",
  1276 => x"0d047198",
  1277 => x"0c04ffb0",
  1278 => x"08b7ec0c",
  1279 => x"04810bff",
  1280 => x"b00c0480",
  1281 => x"0bffb00c",
  1282 => x"0402fc05",
  1283 => x"0d800bb7",
  1284 => x"e80c8051",
  1285 => x"84e52d02",
  1286 => x"84050d04",
  1287 => x"02ec050d",
  1288 => x"76548052",
  1289 => x"870b8815",
  1290 => x"80f52d56",
  1291 => x"53747224",
  1292 => x"8338a053",
  1293 => x"725182ee",
  1294 => x"2d81128b",
  1295 => x"1580f52d",
  1296 => x"54527272",
  1297 => x"25de3802",
  1298 => x"94050d04",
  1299 => x"02f0050d",
  1300 => x"bd980854",
  1301 => x"81f72d80",
  1302 => x"0bbd9c0c",
  1303 => x"7308802e",
  1304 => x"81803882",
  1305 => x"0bb8800c",
  1306 => x"bd9c088f",
  1307 => x"06b7fc0c",
  1308 => x"73085271",
  1309 => x"832e9638",
  1310 => x"71832689",
  1311 => x"3871812e",
  1312 => x"af38a9cd",
  1313 => x"0471852e",
  1314 => x"9f38a9cd",
  1315 => x"04881480",
  1316 => x"f52d8415",
  1317 => x"08b4c053",
  1318 => x"545285f3",
  1319 => x"2d718429",
  1320 => x"13700852",
  1321 => x"52a9d104",
  1322 => x"7351a89c",
  1323 => x"2da9cd04",
  1324 => x"bd940888",
  1325 => x"15082c70",
  1326 => x"81065152",
  1327 => x"71802e87",
  1328 => x"38b4c451",
  1329 => x"a9ca04b4",
  1330 => x"c85185f3",
  1331 => x"2d841408",
  1332 => x"5185f32d",
  1333 => x"bd9c0881",
  1334 => x"05bd9c0c",
  1335 => x"8c1454a8",
  1336 => x"dc040290",
  1337 => x"050d0471",
  1338 => x"bd980ca8",
  1339 => x"cc2dbd9c",
  1340 => x"08ff05bd",
  1341 => x"a00c0402",
  1342 => x"ec050dbd",
  1343 => x"98085580",
  1344 => x"f851a7b9",
  1345 => x"2db7ec08",
  1346 => x"812a7081",
  1347 => x"06515271",
  1348 => x"9b388751",
  1349 => x"a7b92db7",
  1350 => x"ec08812a",
  1351 => x"70810651",
  1352 => x"5271802e",
  1353 => x"b138aaac",
  1354 => x"04a6822d",
  1355 => x"8751a7b9",
  1356 => x"2db7ec08",
  1357 => x"f438aabc",
  1358 => x"04a6822d",
  1359 => x"80f851a7",
  1360 => x"b92db7ec",
  1361 => x"08f338b7",
  1362 => x"e8088132",
  1363 => x"70b7e80c",
  1364 => x"70525284",
  1365 => x"e52db7e8",
  1366 => x"08a23880",
  1367 => x"da51a7b9",
  1368 => x"2d81f551",
  1369 => x"a7b92d81",
  1370 => x"f251a7b9",
  1371 => x"2d81eb51",
  1372 => x"a7b92d81",
  1373 => x"f451a7b9",
  1374 => x"2daec004",
  1375 => x"81f551a7",
  1376 => x"b92db7ec",
  1377 => x"08812a70",
  1378 => x"81065152",
  1379 => x"71802e8f",
  1380 => x"38bda008",
  1381 => x"5271802e",
  1382 => x"8638ff12",
  1383 => x"bda00c81",
  1384 => x"f251a7b9",
  1385 => x"2db7ec08",
  1386 => x"812a7081",
  1387 => x"06515271",
  1388 => x"802e9538",
  1389 => x"bd9c08ff",
  1390 => x"05bda008",
  1391 => x"54527272",
  1392 => x"25863881",
  1393 => x"13bda00c",
  1394 => x"bda00870",
  1395 => x"53547380",
  1396 => x"2e8a388c",
  1397 => x"15ff1555",
  1398 => x"55abce04",
  1399 => x"820bb880",
  1400 => x"0c718f06",
  1401 => x"b7fc0c81",
  1402 => x"eb51a7b9",
  1403 => x"2db7ec08",
  1404 => x"812a7081",
  1405 => x"06515271",
  1406 => x"802ead38",
  1407 => x"7408852e",
  1408 => x"098106a4",
  1409 => x"38881580",
  1410 => x"f52dff05",
  1411 => x"52718816",
  1412 => x"81b72d71",
  1413 => x"982b5271",
  1414 => x"80258838",
  1415 => x"800b8816",
  1416 => x"81b72d74",
  1417 => x"51a89c2d",
  1418 => x"81f451a7",
  1419 => x"b92db7ec",
  1420 => x"08812a70",
  1421 => x"81065152",
  1422 => x"71802eb3",
  1423 => x"38740885",
  1424 => x"2e098106",
  1425 => x"aa388815",
  1426 => x"80f52d81",
  1427 => x"05527188",
  1428 => x"1681b72d",
  1429 => x"7181ff06",
  1430 => x"8b1680f5",
  1431 => x"2d545272",
  1432 => x"72278738",
  1433 => x"72881681",
  1434 => x"b72d7451",
  1435 => x"a89c2d80",
  1436 => x"da51a7b9",
  1437 => x"2db7ec08",
  1438 => x"812a7081",
  1439 => x"06515271",
  1440 => x"802e80fb",
  1441 => x"38bd9808",
  1442 => x"bda00855",
  1443 => x"5373802e",
  1444 => x"8a388c13",
  1445 => x"ff155553",
  1446 => x"ad8d0472",
  1447 => x"08527182",
  1448 => x"2ea63871",
  1449 => x"82268938",
  1450 => x"71812ea5",
  1451 => x"38adff04",
  1452 => x"71832ead",
  1453 => x"3871842e",
  1454 => x"09810680",
  1455 => x"c2388813",
  1456 => x"0851a9e7",
  1457 => x"2dadff04",
  1458 => x"88130852",
  1459 => x"712dadff",
  1460 => x"04810b88",
  1461 => x"14082bbd",
  1462 => x"940832bd",
  1463 => x"940cadfc",
  1464 => x"04881380",
  1465 => x"f52d8105",
  1466 => x"8b1480f5",
  1467 => x"2d535471",
  1468 => x"74248338",
  1469 => x"80547388",
  1470 => x"1481b72d",
  1471 => x"a8cc2d80",
  1472 => x"54800bb8",
  1473 => x"800c738f",
  1474 => x"06b7fc0c",
  1475 => x"a05273bd",
  1476 => x"a0082e09",
  1477 => x"81069838",
  1478 => x"bd9c08ff",
  1479 => x"05743270",
  1480 => x"09810570",
  1481 => x"72079f2a",
  1482 => x"91713151",
  1483 => x"51535371",
  1484 => x"5182ee2d",
  1485 => x"8114548e",
  1486 => x"7425c638",
  1487 => x"b7e80852",
  1488 => x"71b7ec0c",
  1489 => x"0294050d",
  1490 => x"04000000",
  1491 => x"00ffffff",
  1492 => x"ff00ffff",
  1493 => x"ffff00ff",
  1494 => x"ffffff00",
  1495 => x"52657365",
  1496 => x"74000000",
  1497 => x"53617665",
  1498 => x"20616e64",
  1499 => x"20526573",
  1500 => x"65740000",
  1501 => x"4f707469",
  1502 => x"6f6e7320",
  1503 => x"10000000",
  1504 => x"536f756e",
  1505 => x"64201000",
  1506 => x"54757262",
  1507 => x"6f000000",
  1508 => x"4d6f7573",
  1509 => x"6520656d",
  1510 => x"756c6174",
  1511 => x"696f6e00",
  1512 => x"45786974",
  1513 => x"00000000",
  1514 => x"4d617374",
  1515 => x"65720000",
  1516 => x"4f504c4c",
  1517 => x"00000000",
  1518 => x"53434300",
  1519 => x"50534700",
  1520 => x"4261636b",
  1521 => x"00000000",
  1522 => x"5363616e",
  1523 => x"6c696e65",
  1524 => x"73000000",
  1525 => x"53442043",
  1526 => x"61726400",
  1527 => x"4a617061",
  1528 => x"6e657365",
  1529 => x"206b6579",
  1530 => x"206c6179",
  1531 => x"6f757400",
  1532 => x"32303438",
  1533 => x"4c422052",
  1534 => x"414d0000",
  1535 => x"34303936",
  1536 => x"4b422052",
  1537 => x"414d0000",
  1538 => x"536c323a",
  1539 => x"204e6f6e",
  1540 => x"65000000",
  1541 => x"536c323a",
  1542 => x"20455345",
  1543 => x"2d534343",
  1544 => x"20314d42",
  1545 => x"2f534343",
  1546 => x"2d490000",
  1547 => x"536c323a",
  1548 => x"20455345",
  1549 => x"2d52414d",
  1550 => x"20314d42",
  1551 => x"2f415343",
  1552 => x"49493800",
  1553 => x"536c323a",
  1554 => x"20455345",
  1555 => x"2d52414d",
  1556 => x"20314d42",
  1557 => x"2f415343",
  1558 => x"49493136",
  1559 => x"00000000",
  1560 => x"536c313a",
  1561 => x"204e6f6e",
  1562 => x"65000000",
  1563 => x"536c313a",
  1564 => x"20455345",
  1565 => x"2d534343",
  1566 => x"20314d42",
  1567 => x"2f534343",
  1568 => x"2d490000",
  1569 => x"536c313a",
  1570 => x"204d6567",
  1571 => x"6152414d",
  1572 => x"00000000",
  1573 => x"56474120",
  1574 => x"2d203331",
  1575 => x"4b487a2c",
  1576 => x"20363048",
  1577 => x"7a000000",
  1578 => x"56474120",
  1579 => x"2d203331",
  1580 => x"4b487a2c",
  1581 => x"20353048",
  1582 => x"7a000000",
  1583 => x"5456202d",
  1584 => x"20343830",
  1585 => x"692c2036",
  1586 => x"30487a00",
  1587 => x"496e6974",
  1588 => x"69616c69",
  1589 => x"7a696e67",
  1590 => x"20534420",
  1591 => x"63617264",
  1592 => x"0a000000",
  1593 => x"53444843",
  1594 => x"206e6f74",
  1595 => x"20737570",
  1596 => x"706f7274",
  1597 => x"65643b00",
  1598 => x"46617433",
  1599 => x"32206e6f",
  1600 => x"74207375",
  1601 => x"70706f72",
  1602 => x"7465643b",
  1603 => x"00000000",
  1604 => x"0a646973",
  1605 => x"61626c69",
  1606 => x"6e672053",
  1607 => x"44206361",
  1608 => x"72640a10",
  1609 => x"204f4b0a",
  1610 => x"00000000",
  1611 => x"4f434d53",
  1612 => x"58202020",
  1613 => x"43464700",
  1614 => x"54727969",
  1615 => x"6e67204d",
  1616 => x"53583342",
  1617 => x"494f532e",
  1618 => x"5359530a",
  1619 => x"00000000",
  1620 => x"4d535833",
  1621 => x"42494f53",
  1622 => x"53595300",
  1623 => x"54727969",
  1624 => x"6e672042",
  1625 => x"494f535f",
  1626 => x"4d32502e",
  1627 => x"524f4d0a",
  1628 => x"00000000",
  1629 => x"42494f53",
  1630 => x"5f4d3250",
  1631 => x"524f4d00",
  1632 => x"4c6f6164",
  1633 => x"696e6720",
  1634 => x"42494f53",
  1635 => x"0a000000",
  1636 => x"52656164",
  1637 => x"20666169",
  1638 => x"6c65640a",
  1639 => x"00000000",
  1640 => x"4c6f6164",
  1641 => x"696e6720",
  1642 => x"42494f53",
  1643 => x"20666169",
  1644 => x"6c65640a",
  1645 => x"00000000",
  1646 => x"4d425220",
  1647 => x"6661696c",
  1648 => x"0a000000",
  1649 => x"46415431",
  1650 => x"36202020",
  1651 => x"00000000",
  1652 => x"46415433",
  1653 => x"32202020",
  1654 => x"00000000",
  1655 => x"4e6f2070",
  1656 => x"61727469",
  1657 => x"74696f6e",
  1658 => x"20736967",
  1659 => x"0a000000",
  1660 => x"42616420",
  1661 => x"70617274",
  1662 => x"0a000000",
  1663 => x"53444843",
  1664 => x"20657272",
  1665 => x"6f72210a",
  1666 => x"00000000",
  1667 => x"53442069",
  1668 => x"6e69742e",
  1669 => x"2e2e0a00",
  1670 => x"53442063",
  1671 => x"61726420",
  1672 => x"72657365",
  1673 => x"74206661",
  1674 => x"696c6564",
  1675 => x"210a0000",
  1676 => x"57726974",
  1677 => x"65206661",
  1678 => x"696c6564",
  1679 => x"0a000000",
  1680 => x"16200000",
  1681 => x"14200000",
  1682 => x"15200000",
  1683 => x"00000002",
  1684 => x"00000002",
  1685 => x"0000175c",
  1686 => x"0000067f",
  1687 => x"00000002",
  1688 => x"00001764",
  1689 => x"00000671",
  1690 => x"00000004",
  1691 => x"00001774",
  1692 => x"00001af8",
  1693 => x"00000004",
  1694 => x"00001780",
  1695 => x"00001ab0",
  1696 => x"00000001",
  1697 => x"00001788",
  1698 => x"00000007",
  1699 => x"00000001",
  1700 => x"00001790",
  1701 => x"0000000a",
  1702 => x"00000002",
  1703 => x"000017a0",
  1704 => x"00001409",
  1705 => x"00000000",
  1706 => x"00000000",
  1707 => x"00000000",
  1708 => x"00000005",
  1709 => x"000017a8",
  1710 => x"00000007",
  1711 => x"00000005",
  1712 => x"000017b0",
  1713 => x"00000007",
  1714 => x"00000005",
  1715 => x"000017b8",
  1716 => x"00000007",
  1717 => x"00000005",
  1718 => x"000017bc",
  1719 => x"00000007",
  1720 => x"00000004",
  1721 => x"000017c0",
  1722 => x"00001a50",
  1723 => x"00000000",
  1724 => x"00000000",
  1725 => x"00000000",
  1726 => x"00000003",
  1727 => x"00001b88",
  1728 => x"00000003",
  1729 => x"00000001",
  1730 => x"000017c8",
  1731 => x"0000000b",
  1732 => x"00000001",
  1733 => x"000017d4",
  1734 => x"00000002",
  1735 => x"00000003",
  1736 => x"00001b7c",
  1737 => x"00000003",
  1738 => x"00000003",
  1739 => x"00001b6c",
  1740 => x"00000004",
  1741 => x"00000001",
  1742 => x"000017dc",
  1743 => x"00000006",
  1744 => x"00000003",
  1745 => x"00001b64",
  1746 => x"00000002",
  1747 => x"00000004",
  1748 => x"000017c0",
  1749 => x"00001a50",
  1750 => x"00000000",
  1751 => x"00000000",
  1752 => x"00000000",
  1753 => x"000017f0",
  1754 => x"000017fc",
  1755 => x"00001808",
  1756 => x"00001814",
  1757 => x"0000182c",
  1758 => x"00001844",
  1759 => x"00001860",
  1760 => x"0000186c",
  1761 => x"00001884",
  1762 => x"00001894",
  1763 => x"000018a8",
  1764 => x"000018bc",
  1765 => x"00000003",
  1766 => x"00000000",
  1767 => x"00000000",
  1768 => x"00000000",
  1769 => x"00000000",
  1770 => x"00000000",
  1771 => x"00000000",
  1772 => x"00000000",
  1773 => x"00000000",
  1774 => x"00000000",
  1775 => x"00000000",
  1776 => x"00000000",
  1777 => x"00000000",
  1778 => x"00000000",
  1779 => x"00000000",
  1780 => x"00000000",
  1781 => x"00000000",
  1782 => x"00000000",
  1783 => x"00000000",
  1784 => x"00000000",
  1785 => x"00000000",
  1786 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

