-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b88",
     1 => x"e5040000",
     2 => x"00000000",
     3 => x"00000000",
     4 => x"00000000",
     5 => x"00000000",
     6 => x"00000000",
     7 => x"00000000",
     8 => x"88088c08",
     9 => x"90080b0b",
    10 => x"0b88e108",
    11 => x"2d900c8c",
    12 => x"0c880c04",
    13 => x"00000000",
    14 => x"00000000",
    15 => x"00000000",
    16 => x"71fd0608",
    17 => x"72830609",
    18 => x"81058205",
    19 => x"832b2a83",
    20 => x"ffff0652",
    21 => x"04000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"83ffff73",
    26 => x"83060981",
    27 => x"05820583",
    28 => x"2b2b0906",
    29 => x"7383ffff",
    30 => x"0b0b0b0b",
    31 => x"83a50400",
    32 => x"72098105",
    33 => x"72057373",
    34 => x"09060906",
    35 => x"73097306",
    36 => x"070a8106",
    37 => x"53510400",
    38 => x"00000000",
    39 => x"00000000",
    40 => x"72722473",
    41 => x"732e0753",
    42 => x"51040000",
    43 => x"00000000",
    44 => x"00000000",
    45 => x"00000000",
    46 => x"00000000",
    47 => x"00000000",
    48 => x"71737109",
    49 => x"71068106",
    50 => x"09810572",
    51 => x"0a100a72",
    52 => x"0a100a31",
    53 => x"050a8106",
    54 => x"51515351",
    55 => x"04000000",
    56 => x"72722673",
    57 => x"732e0753",
    58 => x"51040000",
    59 => x"00000000",
    60 => x"00000000",
    61 => x"00000000",
    62 => x"00000000",
    63 => x"00000000",
    64 => x"00000000",
    65 => x"00000000",
    66 => x"00000000",
    67 => x"00000000",
    68 => x"00000000",
    69 => x"00000000",
    70 => x"00000000",
    71 => x"00000000",
    72 => x"0b0b0b88",
    73 => x"ba040000",
    74 => x"00000000",
    75 => x"00000000",
    76 => x"00000000",
    77 => x"00000000",
    78 => x"00000000",
    79 => x"00000000",
    80 => x"720a722b",
    81 => x"0a535104",
    82 => x"00000000",
    83 => x"00000000",
    84 => x"00000000",
    85 => x"00000000",
    86 => x"00000000",
    87 => x"00000000",
    88 => x"72729f06",
    89 => x"0981050b",
    90 => x"0b0b889f",
    91 => x"05040000",
    92 => x"00000000",
    93 => x"00000000",
    94 => x"00000000",
    95 => x"00000000",
    96 => x"72722aff",
    97 => x"739f062a",
    98 => x"0974090a",
    99 => x"8106ff05",
   100 => x"06075351",
   101 => x"04000000",
   102 => x"00000000",
   103 => x"00000000",
   104 => x"71715351",
   105 => x"04067383",
   106 => x"06098105",
   107 => x"8205832b",
   108 => x"0b2b0772",
   109 => x"fc060c51",
   110 => x"51040000",
   111 => x"00000000",
   112 => x"72098105",
   113 => x"72050970",
   114 => x"81050906",
   115 => x"0a810653",
   116 => x"51040000",
   117 => x"00000000",
   118 => x"00000000",
   119 => x"00000000",
   120 => x"72098105",
   121 => x"72050970",
   122 => x"81050906",
   123 => x"0a098106",
   124 => x"53510400",
   125 => x"00000000",
   126 => x"00000000",
   127 => x"00000000",
   128 => x"71098105",
   129 => x"52040000",
   130 => x"00000000",
   131 => x"00000000",
   132 => x"00000000",
   133 => x"00000000",
   134 => x"00000000",
   135 => x"00000000",
   136 => x"72720981",
   137 => x"05055351",
   138 => x"04000000",
   139 => x"00000000",
   140 => x"00000000",
   141 => x"00000000",
   142 => x"00000000",
   143 => x"00000000",
   144 => x"72097206",
   145 => x"73730906",
   146 => x"07535104",
   147 => x"00000000",
   148 => x"00000000",
   149 => x"00000000",
   150 => x"00000000",
   151 => x"00000000",
   152 => x"71fc0608",
   153 => x"72830609",
   154 => x"81058305",
   155 => x"1010102a",
   156 => x"81ff0652",
   157 => x"04000000",
   158 => x"00000000",
   159 => x"00000000",
   160 => x"71fc0608",
   161 => x"0b0b0ba3",
   162 => x"f8738306",
   163 => x"10100508",
   164 => x"060b0b0b",
   165 => x"88a20400",
   166 => x"00000000",
   167 => x"00000000",
   168 => x"88088c08",
   169 => x"90087575",
   170 => x"0b0b0b9f",
   171 => x"982d5050",
   172 => x"88085690",
   173 => x"0c8c0c88",
   174 => x"0c510400",
   175 => x"00000000",
   176 => x"88088c08",
   177 => x"90087575",
   178 => x"0b0b0ba0",
   179 => x"ca2d5050",
   180 => x"88085690",
   181 => x"0c8c0c88",
   182 => x"0c510400",
   183 => x"00000000",
   184 => x"72097081",
   185 => x"0509060a",
   186 => x"8106ff05",
   187 => x"70547106",
   188 => x"73097274",
   189 => x"05ff0506",
   190 => x"07515151",
   191 => x"04000000",
   192 => x"72097081",
   193 => x"0509060a",
   194 => x"098106ff",
   195 => x"05705471",
   196 => x"06730972",
   197 => x"7405ff05",
   198 => x"06075151",
   199 => x"51040000",
   200 => x"05ff0504",
   201 => x"00000000",
   202 => x"00000000",
   203 => x"00000000",
   204 => x"00000000",
   205 => x"00000000",
   206 => x"00000000",
   207 => x"00000000",
   208 => x"04000000",
   209 => x"00000000",
   210 => x"00000000",
   211 => x"00000000",
   212 => x"00000000",
   213 => x"00000000",
   214 => x"00000000",
   215 => x"00000000",
   216 => x"71810552",
   217 => x"04000000",
   218 => x"00000000",
   219 => x"00000000",
   220 => x"00000000",
   221 => x"00000000",
   222 => x"00000000",
   223 => x"00000000",
   224 => x"00000000",
   225 => x"00000000",
   226 => x"00000000",
   227 => x"00000000",
   228 => x"00000000",
   229 => x"00000000",
   230 => x"00000000",
   231 => x"00000000",
   232 => x"02840572",
   233 => x"10100552",
   234 => x"04000000",
   235 => x"00000000",
   236 => x"00000000",
   237 => x"00000000",
   238 => x"00000000",
   239 => x"00000000",
   240 => x"00000000",
   241 => x"00000000",
   242 => x"00000000",
   243 => x"00000000",
   244 => x"00000000",
   245 => x"00000000",
   246 => x"00000000",
   247 => x"00000000",
   248 => x"717105ff",
   249 => x"05715351",
   250 => x"020d0400",
   251 => x"00000000",
   252 => x"00000000",
   253 => x"00000000",
   254 => x"00000000",
   255 => x"00000000",
   256 => x"10101010",
   257 => x"10101010",
   258 => x"10101010",
   259 => x"10101010",
   260 => x"10101010",
   261 => x"10101010",
   262 => x"10101010",
   263 => x"10101053",
   264 => x"51047381",
   265 => x"ff067383",
   266 => x"06098105",
   267 => x"83051010",
   268 => x"102b0772",
   269 => x"fc060c51",
   270 => x"51047272",
   271 => x"80728106",
   272 => x"ff050972",
   273 => x"06057110",
   274 => x"52720a10",
   275 => x"0a5372ed",
   276 => x"38515153",
   277 => x"51040000",
   278 => x"800488da",
   279 => x"04040000",
   280 => x"00000004",
   281 => x"5da9b070",
   282 => x"bf92278b",
   283 => x"38807170",
   284 => x"8405530c",
   285 => x"88e70488",
   286 => x"da5188fd",
   287 => x"0402f805",
   288 => x"0da48851",
   289 => x"9b952d98",
   290 => x"bf2d8808",
   291 => x"802ea038",
   292 => x"a4a0519b",
   293 => x"952d89fb",
   294 => x"2d0b0b0b",
   295 => x"a9b052a4",
   296 => x"b85192ee",
   297 => x"2d880887",
   298 => x"38a4c451",
   299 => x"9b952da4",
   300 => x"dc519b95",
   301 => x"2d800b88",
   302 => x"0c028805",
   303 => x"0d0402e8",
   304 => x"050d7779",
   305 => x"7b585555",
   306 => x"80537276",
   307 => x"25a33874",
   308 => x"70810556",
   309 => x"84e02d74",
   310 => x"70810556",
   311 => x"84e02d52",
   312 => x"5271712e",
   313 => x"86388151",
   314 => x"89f30481",
   315 => x"135389ca",
   316 => x"04805170",
   317 => x"880c0298",
   318 => x"050d0402",
   319 => x"d8050dff",
   320 => x"0bbee00c",
   321 => x"800bbef4",
   322 => x"0ca4e851",
   323 => x"9b952dba",
   324 => x"cc528051",
   325 => x"99d52d88",
   326 => x"08548808",
   327 => x"8c38a4f8",
   328 => x"519b952d",
   329 => x"73558fc7",
   330 => x"04a58c51",
   331 => x"9b952d80",
   332 => x"56810bba",
   333 => x"c00c8853",
   334 => x"a5a452bb",
   335 => x"825189be",
   336 => x"2d880876",
   337 => x"2e098106",
   338 => x"86388808",
   339 => x"bac00c88",
   340 => x"53a5b052",
   341 => x"bb9e5189",
   342 => x"be2d8808",
   343 => x"86388808",
   344 => x"bac00cba",
   345 => x"c00852a5",
   346 => x"bc519d98",
   347 => x"2dbac008",
   348 => x"802e8184",
   349 => x"38be920b",
   350 => x"84e02dbe",
   351 => x"930b84e0",
   352 => x"2d71982b",
   353 => x"71902b07",
   354 => x"be940b84",
   355 => x"e02d7088",
   356 => x"2b7207be",
   357 => x"950b84e0",
   358 => x"2d7107be",
   359 => x"ca0b84e0",
   360 => x"2dbecb0b",
   361 => x"84e02d71",
   362 => x"882b0753",
   363 => x"5f54525a",
   364 => x"56575573",
   365 => x"81abaa2e",
   366 => x"0981068c",
   367 => x"3875519b",
   368 => x"dc2d8808",
   369 => x"568bd804",
   370 => x"7382d4d5",
   371 => x"2e8a38a5",
   372 => x"d0519b95",
   373 => x"2d8d8904",
   374 => x"7552a5f0",
   375 => x"519d982d",
   376 => x"bacc5275",
   377 => x"5199d52d",
   378 => x"88085588",
   379 => x"08802e83",
   380 => x"d638a688",
   381 => x"519b952d",
   382 => x"a6b0519d",
   383 => x"982d8853",
   384 => x"a5b052bb",
   385 => x"9e5189be",
   386 => x"2d880889",
   387 => x"38810bbe",
   388 => x"f40c8caf",
   389 => x"048853a5",
   390 => x"a452bb82",
   391 => x"5189be2d",
   392 => x"8808802e",
   393 => x"8a38a6c8",
   394 => x"519d982d",
   395 => x"8d8904be",
   396 => x"ca0b84e0",
   397 => x"2d547380",
   398 => x"d52e0981",
   399 => x"0680ca38",
   400 => x"becb0b84",
   401 => x"e02d5473",
   402 => x"81aa2e09",
   403 => x"8106ba38",
   404 => x"800bbacc",
   405 => x"0b84e02d",
   406 => x"56547481",
   407 => x"e92e8338",
   408 => x"81547481",
   409 => x"eb2e8c38",
   410 => x"80557375",
   411 => x"2e098106",
   412 => x"82d538ba",
   413 => x"d70b84e0",
   414 => x"2d59788d",
   415 => x"38bad80b",
   416 => x"84e02d54",
   417 => x"73822e86",
   418 => x"3880558f",
   419 => x"c704bad9",
   420 => x"0b84e02d",
   421 => x"70befc0c",
   422 => x"ff1170be",
   423 => x"f00c5452",
   424 => x"a6e8519d",
   425 => x"982dbada",
   426 => x"0b84e02d",
   427 => x"badb0b84",
   428 => x"e02d5676",
   429 => x"05758280",
   430 => x"290570be",
   431 => x"e40cbadc",
   432 => x"0b84e02d",
   433 => x"70bedc0c",
   434 => x"bef40859",
   435 => x"57587680",
   436 => x"2e81a438",
   437 => x"8853a5b0",
   438 => x"52bb9e51",
   439 => x"89be2d78",
   440 => x"55880881",
   441 => x"e238befc",
   442 => x"0870842b",
   443 => x"becc0c70",
   444 => x"bef80cba",
   445 => x"f10b84e0",
   446 => x"2dbaf00b",
   447 => x"84e02d71",
   448 => x"82802905",
   449 => x"baf20b84",
   450 => x"e02d7084",
   451 => x"80802912",
   452 => x"baf30b84",
   453 => x"e02d7081",
   454 => x"800a2912",
   455 => x"70bac40c",
   456 => x"bedc0871",
   457 => x"29bee408",
   458 => x"0570bf84",
   459 => x"0cbaf90b",
   460 => x"84e02dba",
   461 => x"f80b84e0",
   462 => x"2d718280",
   463 => x"2905bafa",
   464 => x"0b84e02d",
   465 => x"70848080",
   466 => x"2912bafb",
   467 => x"0b84e02d",
   468 => x"70982b81",
   469 => x"f00a0672",
   470 => x"0570bac8",
   471 => x"0cfe117e",
   472 => x"297705be",
   473 => x"ec0c5257",
   474 => x"52575d57",
   475 => x"51525f52",
   476 => x"5c575757",
   477 => x"8fc504ba",
   478 => x"de0b84e0",
   479 => x"2dbadd0b",
   480 => x"84e02d71",
   481 => x"82802905",
   482 => x"70becc0c",
   483 => x"70a02983",
   484 => x"ff057089",
   485 => x"2a70bef8",
   486 => x"0cbae30b",
   487 => x"84e02dba",
   488 => x"e20b84e0",
   489 => x"2d718280",
   490 => x"290570ba",
   491 => x"c40c7b71",
   492 => x"291e70be",
   493 => x"ec0c7dba",
   494 => x"c80c7305",
   495 => x"bf840c55",
   496 => x"5e515155",
   497 => x"55815574",
   498 => x"880c02a8",
   499 => x"050d0402",
   500 => x"ec050d76",
   501 => x"70872c71",
   502 => x"80ff0657",
   503 => x"5553bef4",
   504 => x"088a3872",
   505 => x"882c7381",
   506 => x"ff065654",
   507 => x"73bee008",
   508 => x"2ea438be",
   509 => x"e4081452",
   510 => x"a78c519d",
   511 => x"982dbacc",
   512 => x"52bee408",
   513 => x"145199d5",
   514 => x"2d880853",
   515 => x"8808802e",
   516 => x"b53873be",
   517 => x"e00cbef4",
   518 => x"08802e97",
   519 => x"38748429",
   520 => x"bacc0570",
   521 => x"0852539b",
   522 => x"dc2d8808",
   523 => x"f00a0655",
   524 => x"90c40474",
   525 => x"10bacc05",
   526 => x"7080c02d",
   527 => x"52539c8b",
   528 => x"2d880855",
   529 => x"74537288",
   530 => x"0c029405",
   531 => x"0d0402c8",
   532 => x"050d7f61",
   533 => x"5f5c8057",
   534 => x"ff0bbee0",
   535 => x"0cbac808",
   536 => x"beec0857",
   537 => x"58bef408",
   538 => x"772e8a38",
   539 => x"befc0884",
   540 => x"2b5990fb",
   541 => x"04bef808",
   542 => x"842b5980",
   543 => x"5a797927",
   544 => x"81ab3879",
   545 => x"8f06a018",
   546 => x"58547397",
   547 => x"387552a7",
   548 => x"ac519d98",
   549 => x"2dbacc52",
   550 => x"75518116",
   551 => x"5699d52d",
   552 => x"bacc5780",
   553 => x"7784e02d",
   554 => x"56547474",
   555 => x"2e833881",
   556 => x"547481e5",
   557 => x"2e80f038",
   558 => x"81707506",
   559 => x"555d7380",
   560 => x"2e80e438",
   561 => x"8b1784e0",
   562 => x"2d98065b",
   563 => x"7a80d838",
   564 => x"8b537d52",
   565 => x"765189be",
   566 => x"2d880880",
   567 => x"ca389c17",
   568 => x"08519bdc",
   569 => x"2d880884",
   570 => x"1d0c9a17",
   571 => x"80c02d51",
   572 => x"9c8b2d88",
   573 => x"08880888",
   574 => x"1e0c8808",
   575 => x"5555bef4",
   576 => x"08802e97",
   577 => x"38941780",
   578 => x"c02d519c",
   579 => x"8b2d8808",
   580 => x"902b83ff",
   581 => x"f00a0670",
   582 => x"16515473",
   583 => x"881d0c7a",
   584 => x"7c0c7c54",
   585 => x"92e60481",
   586 => x"1a5a90fd",
   587 => x"04bef408",
   588 => x"802eb138",
   589 => x"77518fcf",
   590 => x"2d880888",
   591 => x"0853a7cc",
   592 => x"52589d98",
   593 => x"2d7780ff",
   594 => x"fffff806",
   595 => x"547380ff",
   596 => x"fffff82e",
   597 => x"8f38fe18",
   598 => x"befc0829",
   599 => x"bf840805",
   600 => x"5690fb04",
   601 => x"80547388",
   602 => x"0c02b805",
   603 => x"0d0402e4",
   604 => x"050d787a",
   605 => x"7154bed0",
   606 => x"53555590",
   607 => x"ce2d8808",
   608 => x"81ff0653",
   609 => x"72802e80",
   610 => x"e238a7e4",
   611 => x"519b952d",
   612 => x"bed40883",
   613 => x"ff05892a",
   614 => x"57807056",
   615 => x"56757725",
   616 => x"80da38be",
   617 => x"d808fe05",
   618 => x"befc0829",
   619 => x"bf840811",
   620 => x"76bef008",
   621 => x"06057554",
   622 => x"525399d5",
   623 => x"2d880880",
   624 => x"2eb43881",
   625 => x"1570bef0",
   626 => x"08065455",
   627 => x"728d38be",
   628 => x"d808518f",
   629 => x"cf2d8808",
   630 => x"bed80c84",
   631 => x"80148117",
   632 => x"57547676",
   633 => x"24ffbc38",
   634 => x"93fc0474",
   635 => x"52a88051",
   636 => x"9d982d93",
   637 => x"fe048808",
   638 => x"5393fe04",
   639 => x"81537288",
   640 => x"0c029c05",
   641 => x"0d0402f4",
   642 => x"050dd452",
   643 => x"81ff720c",
   644 => x"71085381",
   645 => x"ff720c72",
   646 => x"882b83fe",
   647 => x"80067208",
   648 => x"7081ff06",
   649 => x"51525381",
   650 => x"ff720c72",
   651 => x"7107882b",
   652 => x"72087081",
   653 => x"ff065152",
   654 => x"5381ff72",
   655 => x"0c727107",
   656 => x"882b7208",
   657 => x"7081ff06",
   658 => x"7207880c",
   659 => x"5253028c",
   660 => x"050d0402",
   661 => x"f4050d74",
   662 => x"767181ff",
   663 => x"06d40c53",
   664 => x"53bf8808",
   665 => x"85387189",
   666 => x"2b527198",
   667 => x"2ad40c71",
   668 => x"902a7081",
   669 => x"ff06d40c",
   670 => x"5171882a",
   671 => x"7081ff06",
   672 => x"d40c5171",
   673 => x"81ff06d4",
   674 => x"0c72902a",
   675 => x"7081ff06",
   676 => x"d40c51d4",
   677 => x"087081ff",
   678 => x"06515182",
   679 => x"b8bf5270",
   680 => x"81ff2e09",
   681 => x"81069438",
   682 => x"81ff0bd4",
   683 => x"0cd40870",
   684 => x"81ff06ff",
   685 => x"14545151",
   686 => x"71e53870",
   687 => x"880c028c",
   688 => x"050d0402",
   689 => x"fc050d81",
   690 => x"c75181ff",
   691 => x"0bd40cff",
   692 => x"11517080",
   693 => x"25f43802",
   694 => x"84050d04",
   695 => x"02f0050d",
   696 => x"95c32d81",
   697 => x"9c9f5380",
   698 => x"5287fc80",
   699 => x"f75194d3",
   700 => x"2d880854",
   701 => x"8808812e",
   702 => x"098106a2",
   703 => x"3881ff0b",
   704 => x"d40c820a",
   705 => x"52849c80",
   706 => x"e95194d3",
   707 => x"2d88088b",
   708 => x"3881ff0b",
   709 => x"d40c7353",
   710 => x"96a40495",
   711 => x"c32dff13",
   712 => x"5372c438",
   713 => x"72880c02",
   714 => x"90050d04",
   715 => x"02f4050d",
   716 => x"81ff0bd4",
   717 => x"0ca89051",
   718 => x"9b952d93",
   719 => x"53805287",
   720 => x"fc80c151",
   721 => x"94d32d88",
   722 => x"088b3881",
   723 => x"ff0bd40c",
   724 => x"815396de",
   725 => x"0495c32d",
   726 => x"ff135372",
   727 => x"e0387288",
   728 => x"0c028c05",
   729 => x"0d0402f0",
   730 => x"050d95c3",
   731 => x"2d83aa52",
   732 => x"849c80c8",
   733 => x"5194d32d",
   734 => x"88088808",
   735 => x"53a89c52",
   736 => x"539d982d",
   737 => x"72812e09",
   738 => x"81069a38",
   739 => x"94862d88",
   740 => x"0883ffff",
   741 => x"06537283",
   742 => x"aa2ea038",
   743 => x"880852a8",
   744 => x"b4519d98",
   745 => x"2d96ac2d",
   746 => x"97b60481",
   747 => x"5498b704",
   748 => x"a8cc519d",
   749 => x"982d8054",
   750 => x"98b70481",
   751 => x"ff0bd40c",
   752 => x"b15395dc",
   753 => x"2d880880",
   754 => x"2e80dd38",
   755 => x"805287fc",
   756 => x"80fa5194",
   757 => x"d32d8808",
   758 => x"80c53888",
   759 => x"0852a8e8",
   760 => x"519d982d",
   761 => x"81ff0bd4",
   762 => x"0cd40870",
   763 => x"81ff0670",
   764 => x"54a8f453",
   765 => x"51539d98",
   766 => x"2d81ff0b",
   767 => x"d40c81ff",
   768 => x"0bd40c81",
   769 => x"ff0bd40c",
   770 => x"81ff0bd4",
   771 => x"0c72862a",
   772 => x"70810670",
   773 => x"56515372",
   774 => x"802e9c38",
   775 => x"97ab0488",
   776 => x"0852a8e8",
   777 => x"519d982d",
   778 => x"72822eff",
   779 => x"8338ff13",
   780 => x"5372ff8e",
   781 => x"38725473",
   782 => x"880c0290",
   783 => x"050d0402",
   784 => x"f4050d81",
   785 => x"0bbf880c",
   786 => x"d008708f",
   787 => x"2a708106",
   788 => x"51515372",
   789 => x"f33872d0",
   790 => x"0c95c32d",
   791 => x"a984519b",
   792 => x"952dd008",
   793 => x"708f2a70",
   794 => x"81065151",
   795 => x"5372f338",
   796 => x"810bd00c",
   797 => x"87538052",
   798 => x"84d480c0",
   799 => x"5194d32d",
   800 => x"8808812e",
   801 => x"94387282",
   802 => x"2e098106",
   803 => x"86388053",
   804 => x"99c804ff",
   805 => x"135372de",
   806 => x"3896e62d",
   807 => x"8808bf88",
   808 => x"0c815287",
   809 => x"fc80d051",
   810 => x"94d32d81",
   811 => x"ff0bd40c",
   812 => x"d008708f",
   813 => x"2a708106",
   814 => x"51515372",
   815 => x"f33872d0",
   816 => x"0c81ff0b",
   817 => x"d40c8153",
   818 => x"72880c02",
   819 => x"8c050d04",
   820 => x"800b880c",
   821 => x"0402e005",
   822 => x"0d797b57",
   823 => x"57805881",
   824 => x"ff0bd40c",
   825 => x"d008708f",
   826 => x"2a708106",
   827 => x"51515473",
   828 => x"f3388281",
   829 => x"0bd00c81",
   830 => x"ff0bd40c",
   831 => x"765287fc",
   832 => x"80d15194",
   833 => x"d32d80db",
   834 => x"c6df5588",
   835 => x"08802e8f",
   836 => x"38880853",
   837 => x"7652a990",
   838 => x"519d982d",
   839 => x"9aec0481",
   840 => x"ff0bd40c",
   841 => x"d4087081",
   842 => x"ff065154",
   843 => x"7381fe2e",
   844 => x"0981069c",
   845 => x"3880ff54",
   846 => x"94862d88",
   847 => x"08767084",
   848 => x"05580cff",
   849 => x"14547380",
   850 => x"25ee3881",
   851 => x"589ad604",
   852 => x"ff155574",
   853 => x"ca3881ff",
   854 => x"0bd40cd0",
   855 => x"08708f2a",
   856 => x"70810651",
   857 => x"515473f3",
   858 => x"3873d00c",
   859 => x"77880c02",
   860 => x"a0050d04",
   861 => x"02f8050d",
   862 => x"7352c008",
   863 => x"70882a70",
   864 => x"81065151",
   865 => x"5170802e",
   866 => x"f13871c0",
   867 => x"0c71880c",
   868 => x"0288050d",
   869 => x"0402e805",
   870 => x"0d807857",
   871 => x"55757084",
   872 => x"05570853",
   873 => x"80547298",
   874 => x"2a73882b",
   875 => x"54527180",
   876 => x"2ea238c0",
   877 => x"0870882a",
   878 => x"70810651",
   879 => x"51517080",
   880 => x"2ef13871",
   881 => x"c00c8115",
   882 => x"81155555",
   883 => x"837425d6",
   884 => x"3871ca38",
   885 => x"74880c02",
   886 => x"98050d04",
   887 => x"02f4050d",
   888 => x"7470882a",
   889 => x"83fe8006",
   890 => x"7072982a",
   891 => x"0772882b",
   892 => x"87fc8080",
   893 => x"0673982b",
   894 => x"81f00a06",
   895 => x"71730707",
   896 => x"880c5651",
   897 => x"5351028c",
   898 => x"050d0402",
   899 => x"f8050d02",
   900 => x"8e0584e0",
   901 => x"2d74882b",
   902 => x"077083ff",
   903 => x"ff06880c",
   904 => x"51028805",
   905 => x"0d0402f8",
   906 => x"050d7370",
   907 => x"902b7190",
   908 => x"2a07880c",
   909 => x"52028805",
   910 => x"0d0402ec",
   911 => x"050d7653",
   912 => x"80557275",
   913 => x"258b38ad",
   914 => x"519af42d",
   915 => x"72098105",
   916 => x"5372802e",
   917 => x"b5388754",
   918 => x"729c2a73",
   919 => x"842b5452",
   920 => x"71802e83",
   921 => x"38815589",
   922 => x"72258738",
   923 => x"b712529c",
   924 => x"f504b012",
   925 => x"5274802e",
   926 => x"86387151",
   927 => x"9af42dff",
   928 => x"14547380",
   929 => x"25d2389d",
   930 => x"8f04b051",
   931 => x"9af42d80",
   932 => x"0b880c02",
   933 => x"94050d04",
   934 => x"02c0050d",
   935 => x"0280c405",
   936 => x"57807078",
   937 => x"7084055a",
   938 => x"0872415f",
   939 => x"5d587c70",
   940 => x"84055e08",
   941 => x"5a805b79",
   942 => x"982a7a88",
   943 => x"2b5b5675",
   944 => x"8638775f",
   945 => x"9f8f047d",
   946 => x"802e81a1",
   947 => x"38805e75",
   948 => x"80e42e8a",
   949 => x"387580f8",
   950 => x"2e098106",
   951 => x"89387684",
   952 => x"1871085e",
   953 => x"58547580",
   954 => x"e42e9f38",
   955 => x"7580e426",
   956 => x"8a387580",
   957 => x"e32ebd38",
   958 => x"9ebf0475",
   959 => x"80f32ea2",
   960 => x"387580f8",
   961 => x"2e89389e",
   962 => x"bf048a53",
   963 => x"9e910490",
   964 => x"53ba8052",
   965 => x"7b519cba",
   966 => x"2d8808ba",
   967 => x"805a559e",
   968 => x"cf047684",
   969 => x"18710870",
   970 => x"545b5854",
   971 => x"9b952d80",
   972 => x"559ecf04",
   973 => x"76841871",
   974 => x"08585854",
   975 => x"9efa04a5",
   976 => x"519af42d",
   977 => x"75519af4",
   978 => x"2d821858",
   979 => x"9f820474",
   980 => x"ff165654",
   981 => x"807425aa",
   982 => x"38787081",
   983 => x"055a84e0",
   984 => x"2d705256",
   985 => x"9af42d81",
   986 => x"18589ecf",
   987 => x"0475a52e",
   988 => x"09810686",
   989 => x"38815e9f",
   990 => x"82047551",
   991 => x"9af42d81",
   992 => x"1858811b",
   993 => x"5b837b25",
   994 => x"fead3875",
   995 => x"fea0387e",
   996 => x"880c0280",
   997 => x"c0050d04",
   998 => x"94080294",
   999 => x"0cf93d0d",
  1000 => x"800b9408",
  1001 => x"fc050c94",
  1002 => x"08880508",
  1003 => x"8025ab38",
  1004 => x"94088805",
  1005 => x"08309408",
  1006 => x"88050c80",
  1007 => x"0b9408f4",
  1008 => x"050c9408",
  1009 => x"fc050888",
  1010 => x"38810b94",
  1011 => x"08f4050c",
  1012 => x"9408f405",
  1013 => x"089408fc",
  1014 => x"050c9408",
  1015 => x"8c050880",
  1016 => x"25ab3894",
  1017 => x"088c0508",
  1018 => x"3094088c",
  1019 => x"050c800b",
  1020 => x"9408f005",
  1021 => x"0c9408fc",
  1022 => x"05088838",
  1023 => x"810b9408",
  1024 => x"f0050c94",
  1025 => x"08f00508",
  1026 => x"9408fc05",
  1027 => x"0c805394",
  1028 => x"088c0508",
  1029 => x"52940888",
  1030 => x"05085181",
  1031 => x"a73f8808",
  1032 => x"709408f8",
  1033 => x"050c5494",
  1034 => x"08fc0508",
  1035 => x"802e8c38",
  1036 => x"9408f805",
  1037 => x"08309408",
  1038 => x"f8050c94",
  1039 => x"08f80508",
  1040 => x"70880c54",
  1041 => x"893d0d94",
  1042 => x"0c049408",
  1043 => x"02940cfb",
  1044 => x"3d0d800b",
  1045 => x"9408fc05",
  1046 => x"0c940888",
  1047 => x"05088025",
  1048 => x"93389408",
  1049 => x"88050830",
  1050 => x"94088805",
  1051 => x"0c810b94",
  1052 => x"08fc050c",
  1053 => x"94088c05",
  1054 => x"0880258c",
  1055 => x"3894088c",
  1056 => x"05083094",
  1057 => x"088c050c",
  1058 => x"81539408",
  1059 => x"8c050852",
  1060 => x"94088805",
  1061 => x"0851ad3f",
  1062 => x"88087094",
  1063 => x"08f8050c",
  1064 => x"549408fc",
  1065 => x"0508802e",
  1066 => x"8c389408",
  1067 => x"f8050830",
  1068 => x"9408f805",
  1069 => x"0c9408f8",
  1070 => x"05087088",
  1071 => x"0c54873d",
  1072 => x"0d940c04",
  1073 => x"94080294",
  1074 => x"0cfd3d0d",
  1075 => x"810b9408",
  1076 => x"fc050c80",
  1077 => x"0b9408f8",
  1078 => x"050c9408",
  1079 => x"8c050894",
  1080 => x"08880508",
  1081 => x"27ac3894",
  1082 => x"08fc0508",
  1083 => x"802ea338",
  1084 => x"800b9408",
  1085 => x"8c050824",
  1086 => x"99389408",
  1087 => x"8c050810",
  1088 => x"94088c05",
  1089 => x"0c9408fc",
  1090 => x"05081094",
  1091 => x"08fc050c",
  1092 => x"c9399408",
  1093 => x"fc050880",
  1094 => x"2e80c938",
  1095 => x"94088c05",
  1096 => x"08940888",
  1097 => x"050826a1",
  1098 => x"38940888",
  1099 => x"05089408",
  1100 => x"8c050831",
  1101 => x"94088805",
  1102 => x"0c9408f8",
  1103 => x"05089408",
  1104 => x"fc050807",
  1105 => x"9408f805",
  1106 => x"0c9408fc",
  1107 => x"0508812a",
  1108 => x"9408fc05",
  1109 => x"0c94088c",
  1110 => x"0508812a",
  1111 => x"94088c05",
  1112 => x"0cffaf39",
  1113 => x"94089005",
  1114 => x"08802e8f",
  1115 => x"38940888",
  1116 => x"05087094",
  1117 => x"08f4050c",
  1118 => x"518d3994",
  1119 => x"08f80508",
  1120 => x"709408f4",
  1121 => x"050c5194",
  1122 => x"08f40508",
  1123 => x"880c853d",
  1124 => x"0d940c04",
  1125 => x"94080294",
  1126 => x"0cff3d0d",
  1127 => x"800b9408",
  1128 => x"fc050c94",
  1129 => x"08880508",
  1130 => x"8106ff11",
  1131 => x"70097094",
  1132 => x"088c0508",
  1133 => x"069408fc",
  1134 => x"05081194",
  1135 => x"08fc050c",
  1136 => x"94088805",
  1137 => x"08812a94",
  1138 => x"0888050c",
  1139 => x"94088c05",
  1140 => x"08109408",
  1141 => x"8c050c51",
  1142 => x"51515194",
  1143 => x"08880508",
  1144 => x"802e8438",
  1145 => x"ffbd3994",
  1146 => x"08fc0508",
  1147 => x"70880c51",
  1148 => x"833d0d94",
  1149 => x"0c040000",
  1150 => x"00ffffff",
  1151 => x"ff00ffff",
  1152 => x"ffff00ff",
  1153 => x"ffffff00",
  1154 => x"496e6974",
  1155 => x"69616c69",
  1156 => x"7a696e67",
  1157 => x"20534420",
  1158 => x"63617264",
  1159 => x"0a000000",
  1160 => x"48756e74",
  1161 => x"696e6720",
  1162 => x"666f7220",
  1163 => x"70617274",
  1164 => x"6974696f",
  1165 => x"6e0a0000",
  1166 => x"42494f53",
  1167 => x"5f5f5f5f",
  1168 => x"53595300",
  1169 => x"4c6f6164",
  1170 => x"696e6720",
  1171 => x"42494f53",
  1172 => x"20666169",
  1173 => x"6c65640a",
  1174 => x"00000000",
  1175 => x"52657475",
  1176 => x"726e696e",
  1177 => x"670a0000",
  1178 => x"52656164",
  1179 => x"696e6720",
  1180 => x"4d42520a",
  1181 => x"00000000",
  1182 => x"52656164",
  1183 => x"206f6620",
  1184 => x"4d425220",
  1185 => x"6661696c",
  1186 => x"65640a00",
  1187 => x"4d425220",
  1188 => x"73756363",
  1189 => x"65737366",
  1190 => x"756c6c79",
  1191 => x"20726561",
  1192 => x"640a0000",
  1193 => x"46415431",
  1194 => x"36202020",
  1195 => x"00000000",
  1196 => x"46415433",
  1197 => x"32202020",
  1198 => x"00000000",
  1199 => x"50617274",
  1200 => x"6974696f",
  1201 => x"6e636f75",
  1202 => x"6e742025",
  1203 => x"640a0000",
  1204 => x"4e6f2070",
  1205 => x"61727469",
  1206 => x"74696f6e",
  1207 => x"20736967",
  1208 => x"6e617475",
  1209 => x"72652066",
  1210 => x"6f756e64",
  1211 => x"0a000000",
  1212 => x"52656164",
  1213 => x"696e6720",
  1214 => x"626f6f74",
  1215 => x"20736563",
  1216 => x"746f7220",
  1217 => x"25640a00",
  1218 => x"52656164",
  1219 => x"20626f6f",
  1220 => x"74207365",
  1221 => x"63746f72",
  1222 => x"2066726f",
  1223 => x"6d206669",
  1224 => x"72737420",
  1225 => x"70617274",
  1226 => x"6974696f",
  1227 => x"6e0a0000",
  1228 => x"48756e74",
  1229 => x"696e6720",
  1230 => x"666f7220",
  1231 => x"66696c65",
  1232 => x"73797374",
  1233 => x"656d0a00",
  1234 => x"556e7375",
  1235 => x"70706f72",
  1236 => x"74656420",
  1237 => x"70617274",
  1238 => x"6974696f",
  1239 => x"6e207479",
  1240 => x"7065210d",
  1241 => x"00000000",
  1242 => x"436c7573",
  1243 => x"74657220",
  1244 => x"73697a65",
  1245 => x"3a202564",
  1246 => x"2c20436c",
  1247 => x"75737465",
  1248 => x"72206d61",
  1249 => x"736b2c20",
  1250 => x"25640a00",
  1251 => x"47657443",
  1252 => x"6c757374",
  1253 => x"65722072",
  1254 => x"65616469",
  1255 => x"6e672073",
  1256 => x"6563746f",
  1257 => x"72202564",
  1258 => x"0a000000",
  1259 => x"52656164",
  1260 => x"696e6720",
  1261 => x"64697265",
  1262 => x"63746f72",
  1263 => x"79207365",
  1264 => x"63746f72",
  1265 => x"2025640a",
  1266 => x"00000000",
  1267 => x"47657446",
  1268 => x"41544c69",
  1269 => x"6e6b2072",
  1270 => x"65747572",
  1271 => x"6e656420",
  1272 => x"25640a00",
  1273 => x"4f70656e",
  1274 => x"65642066",
  1275 => x"696c652c",
  1276 => x"206c6f61",
  1277 => x"64696e67",
  1278 => x"2e2e2e0a",
  1279 => x"00000000",
  1280 => x"43616e27",
  1281 => x"74206f70",
  1282 => x"656e2025",
  1283 => x"730a0000",
  1284 => x"436d645f",
  1285 => x"696e6974",
  1286 => x"0a000000",
  1287 => x"636d645f",
  1288 => x"434d4438",
  1289 => x"20726573",
  1290 => x"706f6e73",
  1291 => x"653a2025",
  1292 => x"640a0000",
  1293 => x"434d4438",
  1294 => x"5f342072",
  1295 => x"6573706f",
  1296 => x"6e73653a",
  1297 => x"2025640a",
  1298 => x"00000000",
  1299 => x"53444843",
  1300 => x"20496e69",
  1301 => x"7469616c",
  1302 => x"697a6174",
  1303 => x"696f6e20",
  1304 => x"6572726f",
  1305 => x"72210a00",
  1306 => x"434d4435",
  1307 => x"38202564",
  1308 => x"0a202000",
  1309 => x"434d4435",
  1310 => x"385f3220",
  1311 => x"25640a20",
  1312 => x"20000000",
  1313 => x"53504920",
  1314 => x"496e6974",
  1315 => x"28290a00",
  1316 => x"52656164",
  1317 => x"20636f6d",
  1318 => x"6d616e64",
  1319 => x"20666169",
  1320 => x"6c656420",
  1321 => x"61742025",
  1322 => x"64202825",
  1323 => x"64290a00",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

