-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b0bb1",
     9 => x"d4080b0b",
    10 => x"0bb1d808",
    11 => x"0b0b0bb1",
    12 => x"dc080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"b1dc0c0b",
    16 => x"0b0bb1d8",
    17 => x"0c0b0b0b",
    18 => x"b1d40c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0ba898",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"b1d470b7",
    57 => x"b0278b38",
    58 => x"80717084",
    59 => x"05530c81",
    60 => x"e2048c51",
    61 => x"8a960402",
    62 => x"fc050df8",
    63 => x"80518f0b",
    64 => x"b1e40c9f",
    65 => x"0bb1e80c",
    66 => x"a0717081",
    67 => x"055334b1",
    68 => x"e808ff05",
    69 => x"b1e80cb1",
    70 => x"e8088025",
    71 => x"eb38b1e4",
    72 => x"08ff05b1",
    73 => x"e40cb1e4",
    74 => x"088025d7",
    75 => x"38028405",
    76 => x"0d0402f0",
    77 => x"050df880",
    78 => x"53f8a054",
    79 => x"83bf5273",
    80 => x"70810555",
    81 => x"33517073",
    82 => x"70810555",
    83 => x"34ff1252",
    84 => x"718025eb",
    85 => x"38fbc053",
    86 => x"9f52a073",
    87 => x"70810555",
    88 => x"34ff1252",
    89 => x"718025f2",
    90 => x"38029005",
    91 => x"0d0402f4",
    92 => x"050d7453",
    93 => x"8e0bb1e4",
    94 => x"08258f38",
    95 => x"82b22db1",
    96 => x"e408ff05",
    97 => x"b1e40c82",
    98 => x"f404b1e4",
    99 => x"08b1e808",
   100 => x"5351728a",
   101 => x"2e098106",
   102 => x"b7387151",
   103 => x"719f24a0",
   104 => x"38b1e408",
   105 => x"a02911f8",
   106 => x"80115151",
   107 => x"a07134b1",
   108 => x"e8088105",
   109 => x"b1e80cb1",
   110 => x"e808519f",
   111 => x"7125e238",
   112 => x"800bb1e8",
   113 => x"0cb1e408",
   114 => x"8105b1e4",
   115 => x"0c83e404",
   116 => x"70a02912",
   117 => x"f8801151",
   118 => x"51727134",
   119 => x"b1e80881",
   120 => x"05b1e80c",
   121 => x"b1e808a0",
   122 => x"2e098106",
   123 => x"8e38800b",
   124 => x"b1e80cb1",
   125 => x"e4088105",
   126 => x"b1e40c02",
   127 => x"8c050d04",
   128 => x"02e8050d",
   129 => x"77795656",
   130 => x"880bfc16",
   131 => x"77712c8f",
   132 => x"06545254",
   133 => x"80537272",
   134 => x"25953871",
   135 => x"53fbe014",
   136 => x"51877134",
   137 => x"8114ff14",
   138 => x"545472f1",
   139 => x"387153f9",
   140 => x"1576712c",
   141 => x"87065351",
   142 => x"71802e8b",
   143 => x"38fbe014",
   144 => x"51717134",
   145 => x"81145472",
   146 => x"8e249538",
   147 => x"8f733153",
   148 => x"fbe01451",
   149 => x"a0713481",
   150 => x"14ff1454",
   151 => x"5472f138",
   152 => x"0298050d",
   153 => x"0402ec05",
   154 => x"0d800bb1",
   155 => x"f00cf68c",
   156 => x"08f69008",
   157 => x"71882c57",
   158 => x"5481ff06",
   159 => x"52747225",
   160 => x"88387155",
   161 => x"820bb1f0",
   162 => x"0c72882c",
   163 => x"7381ff06",
   164 => x"54547373",
   165 => x"258b3872",
   166 => x"b1f00884",
   167 => x"07b1f00c",
   168 => x"54b1ec08",
   169 => x"82055182",
   170 => x"0bb1ec0c",
   171 => x"830bf688",
   172 => x"0c74712b",
   173 => x"fecc0570",
   174 => x"9f2a1170",
   175 => x"812c7688",
   176 => x"29ff9405",
   177 => x"70812cb1",
   178 => x"f0085257",
   179 => x"52545151",
   180 => x"76802e85",
   181 => x"38708107",
   182 => x"5170f694",
   183 => x"0c710981",
   184 => x"05f6800c",
   185 => x"72098105",
   186 => x"f6840c02",
   187 => x"94050d04",
   188 => x"02f4050d",
   189 => x"74537270",
   190 => x"81055480",
   191 => x"f52d5271",
   192 => x"802e8938",
   193 => x"715182ee",
   194 => x"2d85f604",
   195 => x"028c050d",
   196 => x"0402d405",
   197 => x"0daafc51",
   198 => x"85f02dab",
   199 => x"9452b1f4",
   200 => x"5192d52d",
   201 => x"b1d40881",
   202 => x"ff065372",
   203 => x"9f38aba0",
   204 => x"5185f02d",
   205 => x"abb852b1",
   206 => x"f45192d5",
   207 => x"2db1d408",
   208 => x"81ff0670",
   209 => x"55537280",
   210 => x"2e81ae38",
   211 => x"abc45185",
   212 => x"f02db1f8",
   213 => x"08578077",
   214 => x"595a767a",
   215 => x"2e8b3881",
   216 => x"1a78812a",
   217 => x"595a77f7",
   218 => x"38f71a5a",
   219 => x"80772581",
   220 => x"81387952",
   221 => x"77518480",
   222 => x"2db28052",
   223 => x"b1f45195",
   224 => x"9a2db1d4",
   225 => x"0881ff06",
   226 => x"5372802e",
   227 => x"80c938b2",
   228 => x"805b8059",
   229 => x"87c4047a",
   230 => x"7084055c",
   231 => x"087081ff",
   232 => x"0671882c",
   233 => x"7081ff06",
   234 => x"73902c70",
   235 => x"81ff0675",
   236 => x"982afec8",
   237 => x"0cfec80c",
   238 => x"58fec80c",
   239 => x"57fec80c",
   240 => x"841a5a53",
   241 => x"76538480",
   242 => x"77258438",
   243 => x"84805372",
   244 => x"7924c438",
   245 => x"87e204ab",
   246 => x"e05185f0",
   247 => x"2d725487",
   248 => x"f904b1f4",
   249 => x"5194ed2d",
   250 => x"fc801781",
   251 => x"19595786",
   252 => x"ec04820b",
   253 => x"fec40c81",
   254 => x"5473b1d4",
   255 => x"0c02ac05",
   256 => x"0d0402f8",
   257 => x"050da3f5",
   258 => x"2d81f72d",
   259 => x"815184e5",
   260 => x"2dfec452",
   261 => x"81720ca1",
   262 => x"bb2da1bb",
   263 => x"2d84720c",
   264 => x"86912d0b",
   265 => x"0b0bafb8",
   266 => x"51a58e2d",
   267 => x"805184e5",
   268 => x"2d028805",
   269 => x"0d0402f4",
   270 => x"050d7470",
   271 => x"8432b7a0",
   272 => x"0c708306",
   273 => x"525370af",
   274 => x"e80b8805",
   275 => x"81b72d72",
   276 => x"892a7081",
   277 => x"06515170",
   278 => x"b0b80b81",
   279 => x"b72d7283",
   280 => x"2a810673",
   281 => x"882a7081",
   282 => x"06515252",
   283 => x"70802e85",
   284 => x"38718207",
   285 => x"5271b088",
   286 => x"0b81b72d",
   287 => x"72842c70",
   288 => x"83065151",
   289 => x"70b0940b",
   290 => x"81b72d70",
   291 => x"b1d40c02",
   292 => x"8c050d04",
   293 => x"02f4050d",
   294 => x"b7a00881",
   295 => x"c406b0b8",
   296 => x"0b80f52d",
   297 => x"52527080",
   298 => x"2e863871",
   299 => x"84800752",
   300 => x"aff00b80",
   301 => x"f52d7207",
   302 => x"b0880b80",
   303 => x"f52d7081",
   304 => x"2a708106",
   305 => x"51535452",
   306 => x"70802e86",
   307 => x"38718280",
   308 => x"07527281",
   309 => x"06517080",
   310 => x"2e853871",
   311 => x"880752b0",
   312 => x"940b80f5",
   313 => x"2d70842b",
   314 => x"73078432",
   315 => x"b1d40c51",
   316 => x"028c050d",
   317 => x"0402f805",
   318 => x"0da1ee2d",
   319 => x"80da51a3",
   320 => x"a52db1d4",
   321 => x"08812a70",
   322 => x"81065152",
   323 => x"71802ee9",
   324 => x"38028805",
   325 => x"0d0402f4",
   326 => x"050d810b",
   327 => x"fec40c84",
   328 => x"b90bfec0",
   329 => x"0c840bfe",
   330 => x"c40ca1d6",
   331 => x"2da3e92d",
   332 => x"a1bb2da1",
   333 => x"bb2d81f7",
   334 => x"2d815184",
   335 => x"e52da1bb",
   336 => x"2da1bb2d",
   337 => x"815184e5",
   338 => x"2dabf451",
   339 => x"85f02d99",
   340 => x"f02db1d4",
   341 => x"08802e81",
   342 => x"923884b9",
   343 => x"528cb92d",
   344 => x"b1d40853",
   345 => x"b1d40880",
   346 => x"2e818738",
   347 => x"9cb22db1",
   348 => x"d408802e",
   349 => x"8738ac8c",
   350 => x"518b8904",
   351 => x"95d12db1",
   352 => x"d408802e",
   353 => x"8d38accc",
   354 => x"5185f02d",
   355 => x"89f52d84",
   356 => x"bd52810b",
   357 => x"fec40c71",
   358 => x"5188b62d",
   359 => x"71fec00c",
   360 => x"840bfec4",
   361 => x"0c86912d",
   362 => x"b1d40880",
   363 => x"2eb73880",
   364 => x"5184e52d",
   365 => x"0b0b0baf",
   366 => x"b851a58e",
   367 => x"2da1ee2d",
   368 => x"a59e2db1",
   369 => x"d4085389",
   370 => x"942db1d4",
   371 => x"08fec00c",
   372 => x"72802e89",
   373 => x"388a0bfe",
   374 => x"c40c8bbd",
   375 => x"04820bfe",
   376 => x"c40c8bbd",
   377 => x"04ad9451",
   378 => x"85f02d82",
   379 => x"0bfec40c",
   380 => x"805372b1",
   381 => x"d40c028c",
   382 => x"050d0402",
   383 => x"e8050d77",
   384 => x"797b5855",
   385 => x"55805372",
   386 => x"7625a338",
   387 => x"74708105",
   388 => x"5680f52d",
   389 => x"74708105",
   390 => x"5680f52d",
   391 => x"52527171",
   392 => x"2e863881",
   393 => x"518cb004",
   394 => x"8113538c",
   395 => x"87048051",
   396 => x"70b1d40c",
   397 => x"0298050d",
   398 => x"0402d805",
   399 => x"0d800bb6",
   400 => x"880cb280",
   401 => x"5280519b",
   402 => x"8f2db1d4",
   403 => x"0854b1d4",
   404 => x"088c38ad",
   405 => x"ac5185f0",
   406 => x"2d735591",
   407 => x"de048056",
   408 => x"810bb6ac",
   409 => x"0c8853ad",
   410 => x"c052b2b6",
   411 => x"518bfb2d",
   412 => x"b1d40876",
   413 => x"2e098106",
   414 => x"8738b1d4",
   415 => x"08b6ac0c",
   416 => x"8853adcc",
   417 => x"52b2d251",
   418 => x"8bfb2db1",
   419 => x"d4088738",
   420 => x"b1d408b6",
   421 => x"ac0cb6ac",
   422 => x"0852add8",
   423 => x"519eac2d",
   424 => x"b6ac0880",
   425 => x"2e80f638",
   426 => x"b5c60b80",
   427 => x"f52db5c7",
   428 => x"0b80f52d",
   429 => x"71982b71",
   430 => x"902b07b5",
   431 => x"c80b80f5",
   432 => x"2d70882b",
   433 => x"7207b5c9",
   434 => x"0b80f52d",
   435 => x"7107b5fe",
   436 => x"0b80f52d",
   437 => x"b5ff0b80",
   438 => x"f52d7188",
   439 => x"2b07535f",
   440 => x"54525a56",
   441 => x"57557381",
   442 => x"abaa2e09",
   443 => x"81068d38",
   444 => x"75519d81",
   445 => x"2db1d408",
   446 => x"568e8904",
   447 => x"7382d4d5",
   448 => x"2e8738ad",
   449 => x"f0518eca",
   450 => x"04b28052",
   451 => x"75519b8f",
   452 => x"2db1d408",
   453 => x"55b1d408",
   454 => x"802e83c2",
   455 => x"388853ad",
   456 => x"cc52b2d2",
   457 => x"518bfb2d",
   458 => x"b1d40889",
   459 => x"38810bb6",
   460 => x"880c8ed0",
   461 => x"048853ad",
   462 => x"c052b2b6",
   463 => x"518bfb2d",
   464 => x"b1d40880",
   465 => x"2e8a38ae",
   466 => x"905185f0",
   467 => x"2d8faa04",
   468 => x"b5fe0b80",
   469 => x"f52d5473",
   470 => x"80d52e09",
   471 => x"810680ca",
   472 => x"38b5ff0b",
   473 => x"80f52d54",
   474 => x"7381aa2e",
   475 => x"098106ba",
   476 => x"38800bb2",
   477 => x"800b80f5",
   478 => x"2d565474",
   479 => x"81e92e83",
   480 => x"38815474",
   481 => x"81eb2e8c",
   482 => x"38805573",
   483 => x"752e0981",
   484 => x"0682cb38",
   485 => x"b28b0b80",
   486 => x"f52d5574",
   487 => x"8d38b28c",
   488 => x"0b80f52d",
   489 => x"5473822e",
   490 => x"86388055",
   491 => x"91de04b2",
   492 => x"8d0b80f5",
   493 => x"2d70b680",
   494 => x"0cff05b6",
   495 => x"840cb28e",
   496 => x"0b80f52d",
   497 => x"b28f0b80",
   498 => x"f52d5876",
   499 => x"05778280",
   500 => x"290570b6",
   501 => x"8c0cb290",
   502 => x"0b80f52d",
   503 => x"70b6a00c",
   504 => x"b6880859",
   505 => x"57587680",
   506 => x"2e81a338",
   507 => x"8853adcc",
   508 => x"52b2d251",
   509 => x"8bfb2db1",
   510 => x"d40881e2",
   511 => x"38b68008",
   512 => x"70842bb6",
   513 => x"a40c70b6",
   514 => x"9c0cb2a5",
   515 => x"0b80f52d",
   516 => x"b2a40b80",
   517 => x"f52d7182",
   518 => x"802905b2",
   519 => x"a60b80f5",
   520 => x"2d708480",
   521 => x"802912b2",
   522 => x"a70b80f5",
   523 => x"2d708180",
   524 => x"0a291270",
   525 => x"b6a80cb6",
   526 => x"a0087129",
   527 => x"b68c0805",
   528 => x"70b6900c",
   529 => x"b2ad0b80",
   530 => x"f52db2ac",
   531 => x"0b80f52d",
   532 => x"71828029",
   533 => x"05b2ae0b",
   534 => x"80f52d70",
   535 => x"84808029",
   536 => x"12b2af0b",
   537 => x"80f52d70",
   538 => x"982b81f0",
   539 => x"0a067205",
   540 => x"70b6940c",
   541 => x"fe117e29",
   542 => x"7705b698",
   543 => x"0c525952",
   544 => x"43545e51",
   545 => x"5259525d",
   546 => x"57595791",
   547 => x"dc04b292",
   548 => x"0b80f52d",
   549 => x"b2910b80",
   550 => x"f52d7182",
   551 => x"80290570",
   552 => x"b6a40c70",
   553 => x"a02983ff",
   554 => x"0570892a",
   555 => x"70b69c0c",
   556 => x"b2970b80",
   557 => x"f52db296",
   558 => x"0b80f52d",
   559 => x"71828029",
   560 => x"0570b6a8",
   561 => x"0c7b7129",
   562 => x"1e70b698",
   563 => x"0c7db694",
   564 => x"0c7305b6",
   565 => x"900c555e",
   566 => x"51515555",
   567 => x"815574b1",
   568 => x"d40c02a8",
   569 => x"050d0402",
   570 => x"ec050d76",
   571 => x"70872c71",
   572 => x"80ff0655",
   573 => x"5654b688",
   574 => x"088a3873",
   575 => x"882c7481",
   576 => x"ff065455",
   577 => x"b28052b6",
   578 => x"8c081551",
   579 => x"9b8f2db1",
   580 => x"d40854b1",
   581 => x"d408802e",
   582 => x"b338b688",
   583 => x"08802e98",
   584 => x"38728429",
   585 => x"b2800570",
   586 => x"0852539d",
   587 => x"812db1d4",
   588 => x"08f00a06",
   589 => x"5392ca04",
   590 => x"7210b280",
   591 => x"057080e0",
   592 => x"2d52539d",
   593 => x"b12db1d4",
   594 => x"08537254",
   595 => x"73b1d40c",
   596 => x"0294050d",
   597 => x"0402c805",
   598 => x"0d7f615f",
   599 => x"5b800bb6",
   600 => x"9408b698",
   601 => x"08595d56",
   602 => x"b6880876",
   603 => x"2e8a38b6",
   604 => x"8008842b",
   605 => x"5892fe04",
   606 => x"b69c0884",
   607 => x"2b588059",
   608 => x"78782781",
   609 => x"a938788f",
   610 => x"06a01757",
   611 => x"54738f38",
   612 => x"b2805276",
   613 => x"51811757",
   614 => x"9b8f2db2",
   615 => x"80568076",
   616 => x"80f52d56",
   617 => x"5474742e",
   618 => x"83388154",
   619 => x"7481e52e",
   620 => x"80f63881",
   621 => x"70750655",
   622 => x"5d73802e",
   623 => x"80ea388b",
   624 => x"1680f52d",
   625 => x"98065a79",
   626 => x"80de388b",
   627 => x"537d5275",
   628 => x"518bfb2d",
   629 => x"b1d40880",
   630 => x"cf389c16",
   631 => x"08519d81",
   632 => x"2db1d408",
   633 => x"841c0c9a",
   634 => x"1680e02d",
   635 => x"519db12d",
   636 => x"b1d408b1",
   637 => x"d408881d",
   638 => x"0cb1d408",
   639 => x"5555b688",
   640 => x"08802e98",
   641 => x"38941680",
   642 => x"e02d519d",
   643 => x"b12db1d4",
   644 => x"08902b83",
   645 => x"fff00a06",
   646 => x"70165154",
   647 => x"73881c0c",
   648 => x"797b0c7c",
   649 => x"5494e404",
   650 => x"81195993",
   651 => x"8004b688",
   652 => x"08802eae",
   653 => x"387b5191",
   654 => x"e72db1d4",
   655 => x"08b1d408",
   656 => x"80ffffff",
   657 => x"f806555c",
   658 => x"7380ffff",
   659 => x"fff82e92",
   660 => x"38b1d408",
   661 => x"fe05b680",
   662 => x"0829b690",
   663 => x"08055792",
   664 => x"fe048054",
   665 => x"73b1d40c",
   666 => x"02b8050d",
   667 => x"0402f405",
   668 => x"0d747008",
   669 => x"8105710c",
   670 => x"7008b684",
   671 => x"08065353",
   672 => x"718e3888",
   673 => x"13085191",
   674 => x"e72db1d4",
   675 => x"0888140c",
   676 => x"810bb1d4",
   677 => x"0c028c05",
   678 => x"0d0402f0",
   679 => x"050d7588",
   680 => x"1108fe05",
   681 => x"b6800829",
   682 => x"b6900811",
   683 => x"7208b684",
   684 => x"08060579",
   685 => x"55535454",
   686 => x"9b8f2db1",
   687 => x"d40853b1",
   688 => x"d408802e",
   689 => x"83388153",
   690 => x"72b1d40c",
   691 => x"0290050d",
   692 => x"04b68808",
   693 => x"b1d40c04",
   694 => x"02f4050d",
   695 => x"d45281ff",
   696 => x"720c7108",
   697 => x"5381ff72",
   698 => x"0c72882b",
   699 => x"83fe8006",
   700 => x"72087081",
   701 => x"ff065152",
   702 => x"5381ff72",
   703 => x"0c727107",
   704 => x"882b7208",
   705 => x"7081ff06",
   706 => x"51525381",
   707 => x"ff720c72",
   708 => x"7107882b",
   709 => x"72087081",
   710 => x"ff067207",
   711 => x"b1d40c52",
   712 => x"53028c05",
   713 => x"0d0402f4",
   714 => x"050d7476",
   715 => x"7181ff06",
   716 => x"d40c5353",
   717 => x"b6b00885",
   718 => x"3871892b",
   719 => x"5271982a",
   720 => x"d40c7190",
   721 => x"2a7081ff",
   722 => x"06d40c51",
   723 => x"71882a70",
   724 => x"81ff06d4",
   725 => x"0c517181",
   726 => x"ff06d40c",
   727 => x"72902a70",
   728 => x"81ff06d4",
   729 => x"0c51d408",
   730 => x"7081ff06",
   731 => x"515182b8",
   732 => x"bf527081",
   733 => x"ff2e0981",
   734 => x"06943881",
   735 => x"ff0bd40c",
   736 => x"d4087081",
   737 => x"ff06ff14",
   738 => x"54515171",
   739 => x"e53870b1",
   740 => x"d40c028c",
   741 => x"050d0402",
   742 => x"fc050d81",
   743 => x"c75181ff",
   744 => x"0bd40cff",
   745 => x"11517080",
   746 => x"25f43802",
   747 => x"84050d04",
   748 => x"02f0050d",
   749 => x"97972d81",
   750 => x"9c9f5380",
   751 => x"5287fc80",
   752 => x"f75196a6",
   753 => x"2db1d408",
   754 => x"54b1d408",
   755 => x"812e0981",
   756 => x"06a33881",
   757 => x"ff0bd40c",
   758 => x"820a5284",
   759 => x"9c80e951",
   760 => x"96a62db1",
   761 => x"d4088b38",
   762 => x"81ff0bd4",
   763 => x"0c735397",
   764 => x"fb049797",
   765 => x"2dff1353",
   766 => x"72c13872",
   767 => x"b1d40c02",
   768 => x"90050d04",
   769 => x"02f4050d",
   770 => x"81ff0bd4",
   771 => x"0c935380",
   772 => x"5287fc80",
   773 => x"c15196a6",
   774 => x"2db1d408",
   775 => x"8b3881ff",
   776 => x"0bd40c81",
   777 => x"5398b104",
   778 => x"97972dff",
   779 => x"135372df",
   780 => x"3872b1d4",
   781 => x"0c028c05",
   782 => x"0d0402f0",
   783 => x"050d9797",
   784 => x"2d83aa52",
   785 => x"849c80c8",
   786 => x"5196a62d",
   787 => x"b1d40881",
   788 => x"2e098106",
   789 => x"923895d8",
   790 => x"2db1d408",
   791 => x"83ffff06",
   792 => x"537283aa",
   793 => x"2e973898",
   794 => x"842d98f8",
   795 => x"04815499",
   796 => x"e704aeb0",
   797 => x"5185f02d",
   798 => x"805499e7",
   799 => x"0481ff0b",
   800 => x"d40cb153",
   801 => x"97b02db1",
   802 => x"d408802e",
   803 => x"80ca3880",
   804 => x"5287fc80",
   805 => x"fa5196a6",
   806 => x"2db1d408",
   807 => x"b13881ff",
   808 => x"0bd40cd4",
   809 => x"085381ff",
   810 => x"0bd40c81",
   811 => x"ff0bd40c",
   812 => x"81ff0bd4",
   813 => x"0c81ff0b",
   814 => x"d40c7286",
   815 => x"2a708106",
   816 => x"b1d40856",
   817 => x"51537280",
   818 => x"2e9d3898",
   819 => x"ed04b1d4",
   820 => x"0852aecc",
   821 => x"519eac2d",
   822 => x"72822eff",
   823 => x"9538ff13",
   824 => x"5372ffa0",
   825 => x"38725473",
   826 => x"b1d40c02",
   827 => x"90050d04",
   828 => x"02f4050d",
   829 => x"810bb6b0",
   830 => x"0cd00870",
   831 => x"8f2a7081",
   832 => x"06515153",
   833 => x"72f33872",
   834 => x"d00c9797",
   835 => x"2daed851",
   836 => x"85f02dd0",
   837 => x"08708f2a",
   838 => x"70810651",
   839 => x"515372f3",
   840 => x"38810bd0",
   841 => x"0c875380",
   842 => x"5284d480",
   843 => x"c05196a6",
   844 => x"2db1d408",
   845 => x"812e9a38",
   846 => x"72822e09",
   847 => x"81068c38",
   848 => x"aef45185",
   849 => x"f02d8053",
   850 => x"9b8604ff",
   851 => x"135372d7",
   852 => x"3898ba2d",
   853 => x"b1d408b6",
   854 => x"b00cb1d4",
   855 => x"088b3881",
   856 => x"5287fc80",
   857 => x"d05196a6",
   858 => x"2d81ff0b",
   859 => x"d40cd008",
   860 => x"708f2a70",
   861 => x"81065151",
   862 => x"5372f338",
   863 => x"72d00c81",
   864 => x"ff0bd40c",
   865 => x"815372b1",
   866 => x"d40c028c",
   867 => x"050d0402",
   868 => x"e0050d79",
   869 => x"7b575780",
   870 => x"5881ff0b",
   871 => x"d40cd008",
   872 => x"708f2a70",
   873 => x"81065151",
   874 => x"5473f338",
   875 => x"82810bd0",
   876 => x"0c81ff0b",
   877 => x"d40c7652",
   878 => x"87fc80d1",
   879 => x"5196a62d",
   880 => x"80dbc6df",
   881 => x"55b1d408",
   882 => x"802e9038",
   883 => x"b1d40853",
   884 => x"7652af8c",
   885 => x"519eac2d",
   886 => x"9ca90481",
   887 => x"ff0bd40c",
   888 => x"d4087081",
   889 => x"ff065154",
   890 => x"7381fe2e",
   891 => x"0981069d",
   892 => x"3880ff54",
   893 => x"95d82db1",
   894 => x"d4087670",
   895 => x"8405580c",
   896 => x"ff145473",
   897 => x"8025ed38",
   898 => x"81589c93",
   899 => x"04ff1555",
   900 => x"74c93881",
   901 => x"ff0bd40c",
   902 => x"d008708f",
   903 => x"2a708106",
   904 => x"51515473",
   905 => x"f33873d0",
   906 => x"0c77b1d4",
   907 => x"0c02a005",
   908 => x"0d04b6b0",
   909 => x"08b1d40c",
   910 => x"0402e805",
   911 => x"0d807857",
   912 => x"55757084",
   913 => x"05570853",
   914 => x"80547298",
   915 => x"2a73882b",
   916 => x"54527180",
   917 => x"2ea238c0",
   918 => x"0870882a",
   919 => x"70810651",
   920 => x"51517080",
   921 => x"2ef13871",
   922 => x"c00c8115",
   923 => x"81155555",
   924 => x"837425d6",
   925 => x"3871ca38",
   926 => x"74b1d40c",
   927 => x"0298050d",
   928 => x"0402f405",
   929 => x"0d747088",
   930 => x"2a83fe80",
   931 => x"06707298",
   932 => x"2a077288",
   933 => x"2b87fc80",
   934 => x"80067398",
   935 => x"2b81f00a",
   936 => x"06717307",
   937 => x"07b1d40c",
   938 => x"56515351",
   939 => x"028c050d",
   940 => x"0402f805",
   941 => x"0d028e05",
   942 => x"80f52d74",
   943 => x"882b0770",
   944 => x"83ffff06",
   945 => x"b1d40c51",
   946 => x"0288050d",
   947 => x"0402ec05",
   948 => x"0d765380",
   949 => x"55727525",
   950 => x"8b38ad51",
   951 => x"82ee2d72",
   952 => x"09810553",
   953 => x"72802eb5",
   954 => x"38875472",
   955 => x"9c2a7384",
   956 => x"2b545271",
   957 => x"802e8338",
   958 => x"81558972",
   959 => x"258738b7",
   960 => x"12529e88",
   961 => x"04b01252",
   962 => x"74802e86",
   963 => x"38715182",
   964 => x"ee2dff14",
   965 => x"54738025",
   966 => x"d2389ea2",
   967 => x"04b05182",
   968 => x"ee2d800b",
   969 => x"b1d40c02",
   970 => x"94050d04",
   971 => x"02c0050d",
   972 => x"0280c405",
   973 => x"57807078",
   974 => x"7084055a",
   975 => x"0872415f",
   976 => x"5d587c70",
   977 => x"84055e08",
   978 => x"5a805b79",
   979 => x"982a7a88",
   980 => x"2b5b5675",
   981 => x"8638775f",
   982 => x"a0a4047d",
   983 => x"802e81a2",
   984 => x"38805e75",
   985 => x"80e42e8a",
   986 => x"387580f8",
   987 => x"2e098106",
   988 => x"89387684",
   989 => x"1871085e",
   990 => x"58547580",
   991 => x"e42e9f38",
   992 => x"7580e426",
   993 => x"8a387580",
   994 => x"e32ebe38",
   995 => x"9fd40475",
   996 => x"80f32ea3",
   997 => x"387580f8",
   998 => x"2e89389f",
   999 => x"d4048a53",
  1000 => x"9fa50490",
  1001 => x"53b6b452",
  1002 => x"7b519dcd",
  1003 => x"2db1d408",
  1004 => x"b6b45a55",
  1005 => x"9fe40476",
  1006 => x"84187108",
  1007 => x"70545b58",
  1008 => x"549cb92d",
  1009 => x"80559fe4",
  1010 => x"04768418",
  1011 => x"71085858",
  1012 => x"54a08f04",
  1013 => x"a55182ee",
  1014 => x"2d755182",
  1015 => x"ee2d8218",
  1016 => x"58a09704",
  1017 => x"74ff1656",
  1018 => x"54807425",
  1019 => x"aa387870",
  1020 => x"81055a80",
  1021 => x"f52d7052",
  1022 => x"5682ee2d",
  1023 => x"8118589f",
  1024 => x"e40475a5",
  1025 => x"2e098106",
  1026 => x"8638815e",
  1027 => x"a0970475",
  1028 => x"5182ee2d",
  1029 => x"81185881",
  1030 => x"1b5b837b",
  1031 => x"25feac38",
  1032 => x"75fe9f38",
  1033 => x"7eb1d40c",
  1034 => x"0280c005",
  1035 => x"0d0402fc",
  1036 => x"050d7251",
  1037 => x"80710c80",
  1038 => x"0b84120c",
  1039 => x"0284050d",
  1040 => x"0402f005",
  1041 => x"0d757008",
  1042 => x"84120853",
  1043 => x"5353ff54",
  1044 => x"71712e9b",
  1045 => x"38841308",
  1046 => x"70842914",
  1047 => x"8b1180f5",
  1048 => x"2d841608",
  1049 => x"81118706",
  1050 => x"84180c52",
  1051 => x"56515173",
  1052 => x"b1d40c02",
  1053 => x"90050d04",
  1054 => x"02f8050d",
  1055 => x"a3ef2de0",
  1056 => x"08708b2a",
  1057 => x"70810651",
  1058 => x"52527080",
  1059 => x"2e9d38b6",
  1060 => x"f4087084",
  1061 => x"29b6fc05",
  1062 => x"7381ff06",
  1063 => x"710c5151",
  1064 => x"b6f40881",
  1065 => x"118706b6",
  1066 => x"f40c5180",
  1067 => x"0bb79c0c",
  1068 => x"a3e22da3",
  1069 => x"e92d0288",
  1070 => x"050d0402",
  1071 => x"fc050da3",
  1072 => x"ef2d810b",
  1073 => x"b79c0ca3",
  1074 => x"e92db79c",
  1075 => x"085170fa",
  1076 => x"38028405",
  1077 => x"0d0402fc",
  1078 => x"050db6f4",
  1079 => x"51a0ae2d",
  1080 => x"a0f851a3",
  1081 => x"de2da388",
  1082 => x"2d028405",
  1083 => x"0d0402f4",
  1084 => x"050da2f0",
  1085 => x"04b1d408",
  1086 => x"81f02e09",
  1087 => x"81068938",
  1088 => x"810bb1c8",
  1089 => x"0ca2f004",
  1090 => x"b1d40881",
  1091 => x"e02e0981",
  1092 => x"06893881",
  1093 => x"0bb1cc0c",
  1094 => x"a2f004b1",
  1095 => x"d40852b1",
  1096 => x"cc08802e",
  1097 => x"8838b1d4",
  1098 => x"08818005",
  1099 => x"5271842c",
  1100 => x"728f0653",
  1101 => x"53b1c808",
  1102 => x"802e9938",
  1103 => x"728429b1",
  1104 => x"88057213",
  1105 => x"81712b70",
  1106 => x"09730806",
  1107 => x"730c5153",
  1108 => x"53a2e604",
  1109 => x"728429b1",
  1110 => x"88057213",
  1111 => x"83712b72",
  1112 => x"0807720c",
  1113 => x"5353800b",
  1114 => x"b1cc0c80",
  1115 => x"0bb1c80c",
  1116 => x"b6f451a0",
  1117 => x"c12db1d4",
  1118 => x"08ff24fe",
  1119 => x"f838800b",
  1120 => x"b1d40c02",
  1121 => x"8c050d04",
  1122 => x"02f8050d",
  1123 => x"b188528f",
  1124 => x"51807270",
  1125 => x"8405540c",
  1126 => x"ff115170",
  1127 => x"8025f238",
  1128 => x"0288050d",
  1129 => x"0402f005",
  1130 => x"0d7551a3",
  1131 => x"ef2d7082",
  1132 => x"2cfc06b1",
  1133 => x"88117210",
  1134 => x"9e067108",
  1135 => x"70722a70",
  1136 => x"83068274",
  1137 => x"2b700974",
  1138 => x"06760c54",
  1139 => x"51565753",
  1140 => x"5153a3e9",
  1141 => x"2d71b1d4",
  1142 => x"0c029005",
  1143 => x"0d047198",
  1144 => x"0c04ffb0",
  1145 => x"08b1d40c",
  1146 => x"04810bff",
  1147 => x"b00c0480",
  1148 => x"0bffb00c",
  1149 => x"0402fc05",
  1150 => x"0d800bb1",
  1151 => x"d00c8051",
  1152 => x"84e52d02",
  1153 => x"84050d04",
  1154 => x"02f0050d",
  1155 => x"b7a40854",
  1156 => x"81f72d80",
  1157 => x"0bb7a80c",
  1158 => x"7308802e",
  1159 => x"80eb3882",
  1160 => x"0bb1e80c",
  1161 => x"b7a8088f",
  1162 => x"06b1e40c",
  1163 => x"73085271",
  1164 => x"812ea438",
  1165 => x"71832e09",
  1166 => x"8106b938",
  1167 => x"881480f5",
  1168 => x"2d841508",
  1169 => x"afac5354",
  1170 => x"5285f02d",
  1171 => x"71842913",
  1172 => x"70085252",
  1173 => x"a4f804b7",
  1174 => x"a0088815",
  1175 => x"082c7081",
  1176 => x"06515271",
  1177 => x"802e8738",
  1178 => x"afb051a4",
  1179 => x"f104afb4",
  1180 => x"5185f02d",
  1181 => x"84140851",
  1182 => x"85f02db7",
  1183 => x"a8088105",
  1184 => x"b7a80c8c",
  1185 => x"1454a498",
  1186 => x"04029005",
  1187 => x"0d0471b7",
  1188 => x"a40ca488",
  1189 => x"2db7a808",
  1190 => x"ff05b7ac",
  1191 => x"0c0402f0",
  1192 => x"050d8751",
  1193 => x"a3a52db1",
  1194 => x"d408812a",
  1195 => x"70810651",
  1196 => x"5271802e",
  1197 => x"a038a5bc",
  1198 => x"04a1ee2d",
  1199 => x"8751a3a5",
  1200 => x"2db1d408",
  1201 => x"f438b1d0",
  1202 => x"08813270",
  1203 => x"b1d00c70",
  1204 => x"525284e5",
  1205 => x"2db1d008",
  1206 => x"963880da",
  1207 => x"51a3a52d",
  1208 => x"81f551a3",
  1209 => x"a52d81f2",
  1210 => x"51a3a52d",
  1211 => x"a88c0481",
  1212 => x"f551a3a5",
  1213 => x"2db1d408",
  1214 => x"812a7081",
  1215 => x"06515271",
  1216 => x"802e8f38",
  1217 => x"b7ac0852",
  1218 => x"71802e86",
  1219 => x"38ff12b7",
  1220 => x"ac0c81f2",
  1221 => x"51a3a52d",
  1222 => x"b1d40881",
  1223 => x"2a708106",
  1224 => x"51527180",
  1225 => x"2e9538b7",
  1226 => x"a808ff05",
  1227 => x"b7ac0854",
  1228 => x"52727225",
  1229 => x"86388113",
  1230 => x"b7ac0c80",
  1231 => x"da51a3a5",
  1232 => x"2db1d408",
  1233 => x"812a7081",
  1234 => x"06515271",
  1235 => x"802e80fb",
  1236 => x"38b7a408",
  1237 => x"b7ac0855",
  1238 => x"5373802e",
  1239 => x"8a388c13",
  1240 => x"ff155553",
  1241 => x"a6d90472",
  1242 => x"08527182",
  1243 => x"2ea63871",
  1244 => x"82268938",
  1245 => x"71812ea5",
  1246 => x"38a7cb04",
  1247 => x"71832ead",
  1248 => x"3871842e",
  1249 => x"09810680",
  1250 => x"c2388813",
  1251 => x"0851a58e",
  1252 => x"2da7cb04",
  1253 => x"88130852",
  1254 => x"712da7cb",
  1255 => x"04810b88",
  1256 => x"14082bb7",
  1257 => x"a00832b7",
  1258 => x"a00ca7c8",
  1259 => x"04881380",
  1260 => x"f52d8105",
  1261 => x"8b1480f5",
  1262 => x"2d535471",
  1263 => x"74248338",
  1264 => x"80547388",
  1265 => x"1481b72d",
  1266 => x"a4882d80",
  1267 => x"54800bb1",
  1268 => x"e80c738f",
  1269 => x"06b1e40c",
  1270 => x"a05273b7",
  1271 => x"ac082e09",
  1272 => x"81069838",
  1273 => x"b7a808ff",
  1274 => x"05743270",
  1275 => x"09810570",
  1276 => x"72079f2a",
  1277 => x"91713151",
  1278 => x"51535371",
  1279 => x"5182ee2d",
  1280 => x"8114548e",
  1281 => x"7425c638",
  1282 => x"b1d00852",
  1283 => x"71b1d40c",
  1284 => x"0290050d",
  1285 => x"04000000",
  1286 => x"00ffffff",
  1287 => x"ff00ffff",
  1288 => x"ffff00ff",
  1289 => x"ffffff00",
  1290 => x"44495020",
  1291 => x"53776974",
  1292 => x"63686573",
  1293 => x"20100000",
  1294 => x"52657365",
  1295 => x"74000000",
  1296 => x"45786974",
  1297 => x"00000000",
  1298 => x"53442043",
  1299 => x"61726400",
  1300 => x"4a617061",
  1301 => x"6e657365",
  1302 => x"206b6579",
  1303 => x"626f6172",
  1304 => x"64206c61",
  1305 => x"796f7574",
  1306 => x"00000000",
  1307 => x"54757262",
  1308 => x"6f202831",
  1309 => x"302e3734",
  1310 => x"4d487a29",
  1311 => x"00000000",
  1312 => x"4261636b",
  1313 => x"00000000",
  1314 => x"32303438",
  1315 => x"4c422052",
  1316 => x"414d0000",
  1317 => x"34303936",
  1318 => x"4b422052",
  1319 => x"414d0000",
  1320 => x"536c323a",
  1321 => x"204e6f6e",
  1322 => x"65000000",
  1323 => x"536c323a",
  1324 => x"20455345",
  1325 => x"2d534343",
  1326 => x"20314d42",
  1327 => x"2f534343",
  1328 => x"2d490000",
  1329 => x"536c323a",
  1330 => x"20455345",
  1331 => x"2d52414d",
  1332 => x"20314d42",
  1333 => x"2f415343",
  1334 => x"49493800",
  1335 => x"536c323a",
  1336 => x"20455345",
  1337 => x"2d52414d",
  1338 => x"20314d42",
  1339 => x"2f415343",
  1340 => x"49493136",
  1341 => x"00000000",
  1342 => x"536c313a",
  1343 => x"204e6f6e",
  1344 => x"65000000",
  1345 => x"536c313a",
  1346 => x"20455345",
  1347 => x"2d534343",
  1348 => x"20314d42",
  1349 => x"2f534343",
  1350 => x"2d490000",
  1351 => x"536c313a",
  1352 => x"204d6567",
  1353 => x"6152414d",
  1354 => x"00000000",
  1355 => x"56474120",
  1356 => x"2d203331",
  1357 => x"4b487a2c",
  1358 => x"20363048",
  1359 => x"7a000000",
  1360 => x"56474120",
  1361 => x"2d203331",
  1362 => x"4b487a2c",
  1363 => x"20353048",
  1364 => x"7a000000",
  1365 => x"53434152",
  1366 => x"54202d20",
  1367 => x"31354b48",
  1368 => x"7a2c2035",
  1369 => x"30487a20",
  1370 => x"52474200",
  1371 => x"54562f53",
  1372 => x"6f756e64",
  1373 => x"202d2031",
  1374 => x"35487a00",
  1375 => x"54727969",
  1376 => x"6e67204d",
  1377 => x"53583342",
  1378 => x"494f532e",
  1379 => x"5359532e",
  1380 => x"2e2e0a00",
  1381 => x"4d535833",
  1382 => x"42494f53",
  1383 => x"53595300",
  1384 => x"54727969",
  1385 => x"6e672042",
  1386 => x"494f535f",
  1387 => x"4d32502e",
  1388 => x"524f4d2e",
  1389 => x"2e2e0a00",
  1390 => x"42494f53",
  1391 => x"5f4d3250",
  1392 => x"524f4d00",
  1393 => x"4f70656e",
  1394 => x"65642042",
  1395 => x"494f532c",
  1396 => x"206c6f61",
  1397 => x"64696e67",
  1398 => x"2e2e2e0a",
  1399 => x"00000000",
  1400 => x"52656164",
  1401 => x"20626c6f",
  1402 => x"636b2066",
  1403 => x"61696c65",
  1404 => x"640a0000",
  1405 => x"496e6974",
  1406 => x"69616c69",
  1407 => x"7a696e67",
  1408 => x"20534420",
  1409 => x"63617264",
  1410 => x"0a000000",
  1411 => x"53444843",
  1412 => x"20636172",
  1413 => x"64206465",
  1414 => x"74656374",
  1415 => x"65642062",
  1416 => x"7574206e",
  1417 => x"6f740a73",
  1418 => x"7570706f",
  1419 => x"72746564",
  1420 => x"3b206469",
  1421 => x"7361626c",
  1422 => x"696e6720",
  1423 => x"53442063",
  1424 => x"6172640a",
  1425 => x"10204f4b",
  1426 => x"0a000000",
  1427 => x"46617433",
  1428 => x"32206669",
  1429 => x"6c657379",
  1430 => x"7374656d",
  1431 => x"20646574",
  1432 => x"65637465",
  1433 => x"64206275",
  1434 => x"740a6e6f",
  1435 => x"74207375",
  1436 => x"70706f72",
  1437 => x"7465643b",
  1438 => x"20646973",
  1439 => x"61626c69",
  1440 => x"6e672053",
  1441 => x"44206361",
  1442 => x"72640a10",
  1443 => x"204f4b0a",
  1444 => x"00000000",
  1445 => x"4c6f6164",
  1446 => x"696e6720",
  1447 => x"42494f53",
  1448 => x"20666169",
  1449 => x"6c65640a",
  1450 => x"00000000",
  1451 => x"52656164",
  1452 => x"206f6620",
  1453 => x"4d425220",
  1454 => x"6661696c",
  1455 => x"65640a00",
  1456 => x"46415431",
  1457 => x"36202020",
  1458 => x"00000000",
  1459 => x"46415433",
  1460 => x"32202020",
  1461 => x"00000000",
  1462 => x"25642070",
  1463 => x"61727469",
  1464 => x"74696f6e",
  1465 => x"7320666f",
  1466 => x"756e640a",
  1467 => x"00000000",
  1468 => x"4e6f2070",
  1469 => x"61727469",
  1470 => x"74696f6e",
  1471 => x"20736967",
  1472 => x"6e617475",
  1473 => x"72652066",
  1474 => x"6f756e64",
  1475 => x"0a000000",
  1476 => x"556e7375",
  1477 => x"70706f72",
  1478 => x"74656420",
  1479 => x"70617274",
  1480 => x"6974696f",
  1481 => x"6e207479",
  1482 => x"7065210a",
  1483 => x"00000000",
  1484 => x"53444843",
  1485 => x"20496e69",
  1486 => x"7469616c",
  1487 => x"697a6174",
  1488 => x"696f6e20",
  1489 => x"6572726f",
  1490 => x"72210a00",
  1491 => x"434d4435",
  1492 => x"38202564",
  1493 => x"0a202000",
  1494 => x"496e6974",
  1495 => x"69616c69",
  1496 => x"73696e67",
  1497 => x"20534420",
  1498 => x"63617264",
  1499 => x"2e2e2e0a",
  1500 => x"00000000",
  1501 => x"53442063",
  1502 => x"61726420",
  1503 => x"72657365",
  1504 => x"74206661",
  1505 => x"696c6564",
  1506 => x"210a0000",
  1507 => x"52656164",
  1508 => x"20636f6d",
  1509 => x"6d616e64",
  1510 => x"20666169",
  1511 => x"6c656420",
  1512 => x"61742025",
  1513 => x"64202825",
  1514 => x"64290a00",
  1515 => x"16200000",
  1516 => x"14200000",
  1517 => x"15200000",
  1518 => x"00000004",
  1519 => x"00001428",
  1520 => x"000017e8",
  1521 => x"00000002",
  1522 => x"00001438",
  1523 => x"00000402",
  1524 => x"00000002",
  1525 => x"00001440",
  1526 => x"000011f5",
  1527 => x"00000000",
  1528 => x"00000000",
  1529 => x"00000000",
  1530 => x"00000003",
  1531 => x"00001878",
  1532 => x"00000004",
  1533 => x"00000001",
  1534 => x"00001448",
  1535 => x"00000002",
  1536 => x"00000003",
  1537 => x"0000186c",
  1538 => x"00000003",
  1539 => x"00000003",
  1540 => x"0000185c",
  1541 => x"00000004",
  1542 => x"00000001",
  1543 => x"00001450",
  1544 => x"00000006",
  1545 => x"00000001",
  1546 => x"0000146c",
  1547 => x"00000007",
  1548 => x"00000003",
  1549 => x"00001854",
  1550 => x"00000002",
  1551 => x"00000004",
  1552 => x"00001480",
  1553 => x"000017b8",
  1554 => x"00000000",
  1555 => x"00000000",
  1556 => x"00000000",
  1557 => x"00001488",
  1558 => x"00001494",
  1559 => x"000014a0",
  1560 => x"000014ac",
  1561 => x"000014c4",
  1562 => x"000014dc",
  1563 => x"000014f8",
  1564 => x"00001504",
  1565 => x"0000151c",
  1566 => x"0000152c",
  1567 => x"00001540",
  1568 => x"00001554",
  1569 => x"0000156c",
  1570 => x"00000000",
  1571 => x"00000000",
  1572 => x"00000000",
  1573 => x"00000000",
  1574 => x"00000000",
  1575 => x"00000000",
  1576 => x"00000000",
  1577 => x"00000000",
  1578 => x"00000000",
  1579 => x"00000000",
  1580 => x"00000000",
  1581 => x"00000000",
  1582 => x"00000000",
  1583 => x"00000000",
  1584 => x"00000000",
  1585 => x"00000000",
  1586 => x"00000000",
  1587 => x"00000000",
  1588 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

