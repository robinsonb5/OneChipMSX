-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"80e60400",
     1 => x"00000000",
     2 => x"0b0b0b0b",
     3 => x"84080d80",
     4 => x"04910471",
     5 => x"fd060872",
     6 => x"83060981",
     7 => x"05820583",
     8 => x"2b2a83ff",
     9 => x"ff065204",
    10 => x"71fc0608",
    11 => x"72830609",
    12 => x"81058305",
    13 => x"1010102a",
    14 => x"81ff0652",
    15 => x"0471fc06",
    16 => x"080b0b0b",
    17 => x"98bc7383",
    18 => x"06101005",
    19 => x"08067381",
    20 => x"ff067383",
    21 => x"06098105",
    22 => x"83051010",
    23 => x"102b0772",
    24 => x"fc060c51",
    25 => x"51040284",
    26 => x"050b0b0b",
    27 => x"0b840c91",
    28 => x"0b818c04",
    29 => x"009df470",
    30 => x"a3e6278b",
    31 => x"38807170",
    32 => x"8405530c",
    33 => x"80f70491",
    34 => x"51818c04",
    35 => x"02f8050d",
    36 => x"98cc5193",
    37 => x"c32d90e4",
    38 => x"2d9df408",
    39 => x"802e9f38",
    40 => x"98e45193",
    41 => x"c32d828a",
    42 => x"2d868da0",
    43 => x"5298fc51",
    44 => x"8afd2d9d",
    45 => x"f4088738",
    46 => x"99885193",
    47 => x"c32d99a0",
    48 => x"5193c32d",
    49 => x"800b9df4",
    50 => x"0c028805",
    51 => x"0d0402e8",
    52 => x"050d7779",
    53 => x"7b585555",
    54 => x"80537276",
    55 => x"25a13874",
    56 => x"70810556",
    57 => x"a82d7470",
    58 => x"810556a8",
    59 => x"2d525271",
    60 => x"712e8638",
    61 => x"81518281",
    62 => x"04811353",
    63 => x"81da0480",
    64 => x"51709df4",
    65 => x"0c029805",
    66 => x"0d0402d8",
    67 => x"050dff0b",
    68 => x"a3b40c80",
    69 => x"0ba3c80c",
    70 => x"99ac5193",
    71 => x"c32d9fa0",
    72 => x"52805191",
    73 => x"fe2d9df4",
    74 => x"08549df4",
    75 => x"088c3899",
    76 => x"bc5193c3",
    77 => x"2d735587",
    78 => x"c70499d0",
    79 => x"5193c32d",
    80 => x"8056810b",
    81 => x"9f940c88",
    82 => x"5399e852",
    83 => x"9fd65181",
    84 => x"ce2d9df4",
    85 => x"08762e09",
    86 => x"81068738",
    87 => x"9df4089f",
    88 => x"940c8853",
    89 => x"99f4529f",
    90 => x"f25181ce",
    91 => x"2d9df408",
    92 => x"87389df4",
    93 => x"089f940c",
    94 => x"9f940852",
    95 => x"9a805195",
    96 => x"ca2d9f94",
    97 => x"08802e81",
    98 => x"8138a2e6",
    99 => x"0ba82da2",
   100 => x"e70ba82d",
   101 => x"71982b71",
   102 => x"902b07a2",
   103 => x"e80ba82d",
   104 => x"70882b72",
   105 => x"07a2e90b",
   106 => x"a82d7107",
   107 => x"a39e0ba8",
   108 => x"2da39f0b",
   109 => x"a82d7188",
   110 => x"2b07535f",
   111 => x"54525a56",
   112 => x"57557381",
   113 => x"abaa2e09",
   114 => x"81068d38",
   115 => x"7551948b",
   116 => x"2d9df408",
   117 => x"5683e804",
   118 => x"7382d4d5",
   119 => x"2e8a389a",
   120 => x"945193c3",
   121 => x"2d859804",
   122 => x"75529ab4",
   123 => x"5195ca2d",
   124 => x"9fa05275",
   125 => x"5191fe2d",
   126 => x"9df40855",
   127 => x"9df40880",
   128 => x"2e83c438",
   129 => x"9acc5193",
   130 => x"c32d9af4",
   131 => x"5195ca2d",
   132 => x"885399f4",
   133 => x"529ff251",
   134 => x"81ce2d9d",
   135 => x"f4088938",
   136 => x"810ba3c8",
   137 => x"0c84c304",
   138 => x"885399e8",
   139 => x"529fd651",
   140 => x"81ce2d9d",
   141 => x"f408802e",
   142 => x"8a389b8c",
   143 => x"5195ca2d",
   144 => x"859804a3",
   145 => x"9e0ba82d",
   146 => x"547380d5",
   147 => x"2e098106",
   148 => x"80c638a3",
   149 => x"9f0ba82d",
   150 => x"547381aa",
   151 => x"2e098106",
   152 => x"b738800b",
   153 => x"9fa00ba8",
   154 => x"2d565474",
   155 => x"81e92e83",
   156 => x"38815474",
   157 => x"81eb2e8c",
   158 => x"38805573",
   159 => x"752e0981",
   160 => x"0682c438",
   161 => x"9fab0ba8",
   162 => x"2d59788c",
   163 => x"389fac0b",
   164 => x"a82d5473",
   165 => x"822e8638",
   166 => x"805587c7",
   167 => x"049fad0b",
   168 => x"a82d70a3",
   169 => x"d00cff11",
   170 => x"70a3c40c",
   171 => x"54529bac",
   172 => x"5195ca2d",
   173 => x"9fae0ba8",
   174 => x"2d9faf0b",
   175 => x"a82d5676",
   176 => x"05758280",
   177 => x"290570a3",
   178 => x"b80c9fb0",
   179 => x"0ba82d70",
   180 => x"a3b00ca3",
   181 => x"c8085957",
   182 => x"5876802e",
   183 => x"819d3888",
   184 => x"5399f452",
   185 => x"9ff25181",
   186 => x"ce2d7855",
   187 => x"9df40881",
   188 => x"d638a3d0",
   189 => x"0870842b",
   190 => x"a3a00c70",
   191 => x"a3cc0c9f",
   192 => x"c50ba82d",
   193 => x"9fc40ba8",
   194 => x"2d718280",
   195 => x"29059fc6",
   196 => x"0ba82d70",
   197 => x"84808029",
   198 => x"129fc70b",
   199 => x"a82d7081",
   200 => x"800a2912",
   201 => x"709f980c",
   202 => x"a3b00871",
   203 => x"29a3b808",
   204 => x"0570a3d8",
   205 => x"0c9fcd0b",
   206 => x"a82d9fcc",
   207 => x"0ba82d71",
   208 => x"82802905",
   209 => x"9fce0ba8",
   210 => x"2d708480",
   211 => x"8029129f",
   212 => x"cf0ba82d",
   213 => x"70982b81",
   214 => x"f00a0672",
   215 => x"05709f9c",
   216 => x"0cfe117e",
   217 => x"297705a3",
   218 => x"c00c5257",
   219 => x"52575d57",
   220 => x"51525f52",
   221 => x"5c575757",
   222 => x"87c5049f",
   223 => x"b20ba82d",
   224 => x"9fb10ba8",
   225 => x"2d718280",
   226 => x"290570a3",
   227 => x"a00c70a0",
   228 => x"2983ff05",
   229 => x"70892a70",
   230 => x"a3cc0c9f",
   231 => x"b70ba82d",
   232 => x"9fb60ba8",
   233 => x"2d718280",
   234 => x"2905709f",
   235 => x"980c7b71",
   236 => x"291e70a3",
   237 => x"c00c7d9f",
   238 => x"9c0c7305",
   239 => x"a3d80c55",
   240 => x"5e515155",
   241 => x"55815574",
   242 => x"9df40c02",
   243 => x"a8050d04",
   244 => x"02ec050d",
   245 => x"7670872c",
   246 => x"7180ff06",
   247 => x"575553a3",
   248 => x"c8088a38",
   249 => x"72882c73",
   250 => x"81ff0656",
   251 => x"5473a3b4",
   252 => x"082ea638",
   253 => x"a3b80814",
   254 => x"529bd051",
   255 => x"95ca2d9f",
   256 => x"a052a3b8",
   257 => x"08145191",
   258 => x"fe2d9df4",
   259 => x"08539df4",
   260 => x"08802eb6",
   261 => x"3873a3b4",
   262 => x"0ca3c808",
   263 => x"802e9838",
   264 => x"7484299f",
   265 => x"a0057008",
   266 => x"5253948b",
   267 => x"2d9df408",
   268 => x"f00a0655",
   269 => x"88c80474",
   270 => x"109fa005",
   271 => x"70932d52",
   272 => x"5394bb2d",
   273 => x"9df40855",
   274 => x"7453729d",
   275 => x"f40c0294",
   276 => x"050d0402",
   277 => x"c8050d7f",
   278 => x"615f5c80",
   279 => x"57ff0ba3",
   280 => x"b40c9f9c",
   281 => x"08a3c008",
   282 => x"5758a3c8",
   283 => x"08772e8a",
   284 => x"38a3d008",
   285 => x"842b5989",
   286 => x"8004a3cc",
   287 => x"08842b59",
   288 => x"805a7979",
   289 => x"2781b238",
   290 => x"798f06a0",
   291 => x"18585473",
   292 => x"97387552",
   293 => x"9bf05195",
   294 => x"ca2d9fa0",
   295 => x"52755181",
   296 => x"165691fe",
   297 => x"2d9fa057",
   298 => x"8077a82d",
   299 => x"56547474",
   300 => x"2e833881",
   301 => x"547481e5",
   302 => x"2e80f838",
   303 => x"81707506",
   304 => x"555d7380",
   305 => x"2e80ec38",
   306 => x"8b17a82d",
   307 => x"98065b7a",
   308 => x"80e13876",
   309 => x"5193c32d",
   310 => x"8b537d52",
   311 => x"765181ce",
   312 => x"2d9df408",
   313 => x"80cd389c",
   314 => x"17085194",
   315 => x"8b2d9df4",
   316 => x"08841d0c",
   317 => x"9a17932d",
   318 => x"5194bb2d",
   319 => x"9df4089d",
   320 => x"f408881e",
   321 => x"0c9df408",
   322 => x"5555a3c8",
   323 => x"08802e97",
   324 => x"38941793",
   325 => x"2d5194bb",
   326 => x"2d9df408",
   327 => x"902b83ff",
   328 => x"f00a0670",
   329 => x"16515473",
   330 => x"881d0c7a",
   331 => x"7c0c7c54",
   332 => x"8af40481",
   333 => x"1a5a8982",
   334 => x"04a3c808",
   335 => x"802eb338",
   336 => x"775187d0",
   337 => x"2d9df408",
   338 => x"9df40853",
   339 => x"9c905258",
   340 => x"95ca2d77",
   341 => x"80ffffff",
   342 => x"f8065473",
   343 => x"80ffffff",
   344 => x"f82e8f38",
   345 => x"fe18a3d0",
   346 => x"0829a3d8",
   347 => x"08055689",
   348 => x"80048054",
   349 => x"739df40c",
   350 => x"02b8050d",
   351 => x"0402e405",
   352 => x"0d787a71",
   353 => x"54a3a453",
   354 => x"555588d3",
   355 => x"2d9df408",
   356 => x"81ff0653",
   357 => x"72802e80",
   358 => x"e4389ca8",
   359 => x"5193c32d",
   360 => x"a3a80883",
   361 => x"ff05892a",
   362 => x"57807056",
   363 => x"56757725",
   364 => x"80dd38a3",
   365 => x"ac08fe05",
   366 => x"a3d00829",
   367 => x"a3d80811",
   368 => x"76a3c408",
   369 => x"06057554",
   370 => x"525391fe",
   371 => x"2d9df408",
   372 => x"802eb538",
   373 => x"811570a3",
   374 => x"c4080654",
   375 => x"55728e38",
   376 => x"a3ac0851",
   377 => x"87d02d9d",
   378 => x"f408a3ac",
   379 => x"0c848014",
   380 => x"81175754",
   381 => x"767624ff",
   382 => x"ba388c8f",
   383 => x"0474529c",
   384 => x"c45195ca",
   385 => x"2d8c9104",
   386 => x"9df40853",
   387 => x"8c910481",
   388 => x"53729df4",
   389 => x"0c029c05",
   390 => x"0d0402f4",
   391 => x"050dd452",
   392 => x"81ff720c",
   393 => x"71085381",
   394 => x"ff720c72",
   395 => x"882b83fe",
   396 => x"80067208",
   397 => x"7081ff06",
   398 => x"51525381",
   399 => x"ff720c72",
   400 => x"7107882b",
   401 => x"72087081",
   402 => x"ff065152",
   403 => x"5381ff72",
   404 => x"0c727107",
   405 => x"882b7208",
   406 => x"7081ff06",
   407 => x"72079df4",
   408 => x"0c525302",
   409 => x"8c050d04",
   410 => x"02f4050d",
   411 => x"74767181",
   412 => x"ff06d40c",
   413 => x"5353a3dc",
   414 => x"08853871",
   415 => x"892b5271",
   416 => x"982ad40c",
   417 => x"71902a70",
   418 => x"81ff06d4",
   419 => x"0c517188",
   420 => x"2a7081ff",
   421 => x"06d40c51",
   422 => x"7181ff06",
   423 => x"d40c7290",
   424 => x"2a7081ff",
   425 => x"06d40c51",
   426 => x"d4087081",
   427 => x"ff065151",
   428 => x"82b8bf52",
   429 => x"7081ff2e",
   430 => x"09810694",
   431 => x"3881ff0b",
   432 => x"d40cd408",
   433 => x"7081ff06",
   434 => x"ff145451",
   435 => x"5171e538",
   436 => x"709df40c",
   437 => x"028c050d",
   438 => x"0402fc05",
   439 => x"0d81c751",
   440 => x"81ff0bd4",
   441 => x"0cff1151",
   442 => x"708025f4",
   443 => x"38028405",
   444 => x"0d0402f0",
   445 => x"050d8dd9",
   446 => x"2d819c9f",
   447 => x"53805287",
   448 => x"fc80f751",
   449 => x"8ce82d9d",
   450 => x"f408549d",
   451 => x"f408812e",
   452 => x"098106a3",
   453 => x"3881ff0b",
   454 => x"d40c820a",
   455 => x"52849c80",
   456 => x"e9518ce8",
   457 => x"2d9df408",
   458 => x"8b3881ff",
   459 => x"0bd40c73",
   460 => x"538ebd04",
   461 => x"8dd92dff",
   462 => x"135372c1",
   463 => x"38729df4",
   464 => x"0c029005",
   465 => x"0d0402f4",
   466 => x"050d81ff",
   467 => x"0bd40c9c",
   468 => x"d45193c3",
   469 => x"2d935380",
   470 => x"5287fc80",
   471 => x"c1518ce8",
   472 => x"2d9df408",
   473 => x"8b3881ff",
   474 => x"0bd40c81",
   475 => x"538ef904",
   476 => x"8dd92dff",
   477 => x"135372df",
   478 => x"38729df4",
   479 => x"0c028c05",
   480 => x"0d0402f0",
   481 => x"050d8dd9",
   482 => x"2d83aa52",
   483 => x"849c80c8",
   484 => x"518ce82d",
   485 => x"9df4089d",
   486 => x"f408539c",
   487 => x"e0525395",
   488 => x"ca2d7281",
   489 => x"2e098106",
   490 => x"9c388c9a",
   491 => x"2d9df408",
   492 => x"83ffff06",
   493 => x"537283aa",
   494 => x"2ea1389d",
   495 => x"f408529c",
   496 => x"f85195ca",
   497 => x"2d8ec62d",
   498 => x"8fd60481",
   499 => x"5490db04",
   500 => x"9d905195",
   501 => x"ca2d8054",
   502 => x"90db0481",
   503 => x"ff0bd40c",
   504 => x"b1538df2",
   505 => x"2d9df408",
   506 => x"802e80e0",
   507 => x"38805287",
   508 => x"fc80fa51",
   509 => x"8ce82d9d",
   510 => x"f40880c6",
   511 => x"389df408",
   512 => x"529dac51",
   513 => x"95ca2d81",
   514 => x"ff0bd40c",
   515 => x"d4087081",
   516 => x"ff067054",
   517 => x"9db85351",
   518 => x"5395ca2d",
   519 => x"81ff0bd4",
   520 => x"0c81ff0b",
   521 => x"d40c81ff",
   522 => x"0bd40c81",
   523 => x"ff0bd40c",
   524 => x"72862a70",
   525 => x"81067056",
   526 => x"51537280",
   527 => x"2e9d388f",
   528 => x"cb049df4",
   529 => x"08529dac",
   530 => x"5195ca2d",
   531 => x"72822efe",
   532 => x"ff38ff13",
   533 => x"5372ff8a",
   534 => x"38725473",
   535 => x"9df40c02",
   536 => x"90050d04",
   537 => x"02f4050d",
   538 => x"810ba3dc",
   539 => x"0cd00870",
   540 => x"8f2a7081",
   541 => x"06515153",
   542 => x"72f33872",
   543 => x"d00c8dd9",
   544 => x"2d9dc851",
   545 => x"93c32dd0",
   546 => x"08708f2a",
   547 => x"70810651",
   548 => x"515372f3",
   549 => x"38810bd0",
   550 => x"0c875380",
   551 => x"5284d480",
   552 => x"c0518ce8",
   553 => x"2d9df408",
   554 => x"812e9438",
   555 => x"72822e09",
   556 => x"81068638",
   557 => x"805391ef",
   558 => x"04ff1353",
   559 => x"72dd388f",
   560 => x"822d9df4",
   561 => x"08a3dc0c",
   562 => x"815287fc",
   563 => x"80d0518c",
   564 => x"e82d81ff",
   565 => x"0bd40cd0",
   566 => x"08708f2a",
   567 => x"70810651",
   568 => x"515372f3",
   569 => x"3872d00c",
   570 => x"81ff0bd4",
   571 => x"0c815372",
   572 => x"9df40c02",
   573 => x"8c050d04",
   574 => x"800b9df4",
   575 => x"0c0402e0",
   576 => x"050d797b",
   577 => x"57578058",
   578 => x"81ff0bd4",
   579 => x"0cd00870",
   580 => x"8f2a7081",
   581 => x"06515154",
   582 => x"73f33882",
   583 => x"810bd00c",
   584 => x"81ff0bd4",
   585 => x"0c765287",
   586 => x"fc80d151",
   587 => x"8ce82d80",
   588 => x"dbc6df55",
   589 => x"9df40880",
   590 => x"2e90389d",
   591 => x"f4085376",
   592 => x"529dd451",
   593 => x"95ca2d93",
   594 => x"980481ff",
   595 => x"0bd40cd4",
   596 => x"087081ff",
   597 => x"06515473",
   598 => x"81fe2e09",
   599 => x"81069d38",
   600 => x"80ff548c",
   601 => x"9a2d9df4",
   602 => x"08767084",
   603 => x"05580cff",
   604 => x"14547380",
   605 => x"25ed3881",
   606 => x"58938204",
   607 => x"ff155574",
   608 => x"c93881ff",
   609 => x"0bd40cd0",
   610 => x"08708f2a",
   611 => x"70810651",
   612 => x"515473f3",
   613 => x"3873d00c",
   614 => x"779df40c",
   615 => x"02a0050d",
   616 => x"0402f805",
   617 => x"0d7352c0",
   618 => x"0870882a",
   619 => x"70810651",
   620 => x"51517080",
   621 => x"2ef13871",
   622 => x"c00c719d",
   623 => x"f40c0288",
   624 => x"050d0402",
   625 => x"e8050d80",
   626 => x"78575575",
   627 => x"70840557",
   628 => x"08538054",
   629 => x"72982a73",
   630 => x"882b5452",
   631 => x"71802ea2",
   632 => x"38c00870",
   633 => x"882a7081",
   634 => x"06515151",
   635 => x"70802ef1",
   636 => x"3871c00c",
   637 => x"81158115",
   638 => x"55558374",
   639 => x"25d63871",
   640 => x"ca38749d",
   641 => x"f40c0298",
   642 => x"050d0402",
   643 => x"f4050d74",
   644 => x"70882a83",
   645 => x"fe800670",
   646 => x"72982a07",
   647 => x"72882b87",
   648 => x"fc808006",
   649 => x"73982b81",
   650 => x"f00a0671",
   651 => x"7307079d",
   652 => x"f40c5651",
   653 => x"5351028c",
   654 => x"050d0402",
   655 => x"f8050d02",
   656 => x"8e05a82d",
   657 => x"74882b07",
   658 => x"7083ffff",
   659 => x"069df40c",
   660 => x"51028805",
   661 => x"0d0402f8",
   662 => x"050d7370",
   663 => x"902b7190",
   664 => x"2a079df4",
   665 => x"0c520288",
   666 => x"050d0402",
   667 => x"ec050d76",
   668 => x"53805572",
   669 => x"75258b38",
   670 => x"ad5193a1",
   671 => x"2d720981",
   672 => x"05537280",
   673 => x"2eb53887",
   674 => x"54729c2a",
   675 => x"73842b54",
   676 => x"5271802e",
   677 => x"83388155",
   678 => x"89722587",
   679 => x"38b71252",
   680 => x"95a604b0",
   681 => x"12527480",
   682 => x"2e863871",
   683 => x"5193a12d",
   684 => x"ff145473",
   685 => x"8025d238",
   686 => x"95c004b0",
   687 => x"5193a12d",
   688 => x"800b9df4",
   689 => x"0c029405",
   690 => x"0d0402c0",
   691 => x"050d0280",
   692 => x"c4055780",
   693 => x"70787084",
   694 => x"055a0872",
   695 => x"415f5d58",
   696 => x"7c708405",
   697 => x"5e085a80",
   698 => x"5b79982a",
   699 => x"7a882b5b",
   700 => x"56758638",
   701 => x"775f97c1",
   702 => x"047d802e",
   703 => x"81a13880",
   704 => x"5e7580e4",
   705 => x"2e8a3875",
   706 => x"80f82e09",
   707 => x"81068938",
   708 => x"76841871",
   709 => x"085e5854",
   710 => x"7580e42e",
   711 => x"9f387580",
   712 => x"e4268a38",
   713 => x"7580e32e",
   714 => x"be3896f2",
   715 => x"047580f3",
   716 => x"2ea33875",
   717 => x"80f82e89",
   718 => x"3896f204",
   719 => x"8a5396c3",
   720 => x"0490539e",
   721 => x"d4527b51",
   722 => x"94eb2d9d",
   723 => x"f4089ed4",
   724 => x"5a559782",
   725 => x"04768418",
   726 => x"71087054",
   727 => x"5b585493",
   728 => x"c32d8055",
   729 => x"97820476",
   730 => x"84187108",
   731 => x"58585497",
   732 => x"ac04a551",
   733 => x"93a12d75",
   734 => x"5193a12d",
   735 => x"82185897",
   736 => x"b40474ff",
   737 => x"16565480",
   738 => x"7425a938",
   739 => x"78708105",
   740 => x"5aa82d70",
   741 => x"525693a1",
   742 => x"2d811858",
   743 => x"97820475",
   744 => x"a52e0981",
   745 => x"06863881",
   746 => x"5e97b404",
   747 => x"755193a1",
   748 => x"2d811858",
   749 => x"811b5b83",
   750 => x"7b25fead",
   751 => x"3875fea0",
   752 => x"387e9df4",
   753 => x"0c0280c0",
   754 => x"050d049e",
   755 => x"8008029e",
   756 => x"800cff3d",
   757 => x"0d800b9e",
   758 => x"8008fc05",
   759 => x"0c9e8008",
   760 => x"88050881",
   761 => x"06ff1170",
   762 => x"09709e80",
   763 => x"088c0508",
   764 => x"069e8008",
   765 => x"fc050811",
   766 => x"9e8008fc",
   767 => x"050c9e80",
   768 => x"08880508",
   769 => x"812a9e80",
   770 => x"0888050c",
   771 => x"9e80088c",
   772 => x"0508109e",
   773 => x"80088c05",
   774 => x"0c515151",
   775 => x"519e8008",
   776 => x"88050880",
   777 => x"2e8438ff",
   778 => x"b4399e80",
   779 => x"08fc0508",
   780 => x"709df40c",
   781 => x"51833d0d",
   782 => x"9e800c04",
   783 => x"00ffffff",
   784 => x"ff00ffff",
   785 => x"ffff00ff",
   786 => x"ffffff00",
   787 => x"496e6974",
   788 => x"69616c69",
   789 => x"7a696e67",
   790 => x"20534420",
   791 => x"63617264",
   792 => x"0a000000",
   793 => x"48756e74",
   794 => x"696e6720",
   795 => x"666f7220",
   796 => x"70617274",
   797 => x"6974696f",
   798 => x"6e0a0000",
   799 => x"42494f53",
   800 => x"5f4d3250",
   801 => x"524f4d00",
   802 => x"4c6f6164",
   803 => x"696e6720",
   804 => x"42494f53",
   805 => x"20666169",
   806 => x"6c65640a",
   807 => x"00000000",
   808 => x"52657475",
   809 => x"726e696e",
   810 => x"670a0000",
   811 => x"52656164",
   812 => x"696e6720",
   813 => x"4d42520a",
   814 => x"00000000",
   815 => x"52656164",
   816 => x"206f6620",
   817 => x"4d425220",
   818 => x"6661696c",
   819 => x"65640a00",
   820 => x"4d425220",
   821 => x"73756363",
   822 => x"65737366",
   823 => x"756c6c79",
   824 => x"20726561",
   825 => x"640a0000",
   826 => x"46415431",
   827 => x"36202020",
   828 => x"00000000",
   829 => x"46415433",
   830 => x"32202020",
   831 => x"00000000",
   832 => x"50617274",
   833 => x"6974696f",
   834 => x"6e636f75",
   835 => x"6e742025",
   836 => x"640a0000",
   837 => x"4e6f2070",
   838 => x"61727469",
   839 => x"74696f6e",
   840 => x"20736967",
   841 => x"6e617475",
   842 => x"72652066",
   843 => x"6f756e64",
   844 => x"0a000000",
   845 => x"52656164",
   846 => x"696e6720",
   847 => x"626f6f74",
   848 => x"20736563",
   849 => x"746f7220",
   850 => x"25640a00",
   851 => x"52656164",
   852 => x"20626f6f",
   853 => x"74207365",
   854 => x"63746f72",
   855 => x"2066726f",
   856 => x"6d206669",
   857 => x"72737420",
   858 => x"70617274",
   859 => x"6974696f",
   860 => x"6e0a0000",
   861 => x"48756e74",
   862 => x"696e6720",
   863 => x"666f7220",
   864 => x"66696c65",
   865 => x"73797374",
   866 => x"656d0a00",
   867 => x"556e7375",
   868 => x"70706f72",
   869 => x"74656420",
   870 => x"70617274",
   871 => x"6974696f",
   872 => x"6e207479",
   873 => x"7065210d",
   874 => x"00000000",
   875 => x"436c7573",
   876 => x"74657220",
   877 => x"73697a65",
   878 => x"3a202564",
   879 => x"2c20436c",
   880 => x"75737465",
   881 => x"72206d61",
   882 => x"736b2c20",
   883 => x"25640a00",
   884 => x"47657443",
   885 => x"6c757374",
   886 => x"65722072",
   887 => x"65616469",
   888 => x"6e672073",
   889 => x"6563746f",
   890 => x"72202564",
   891 => x"0a000000",
   892 => x"52656164",
   893 => x"696e6720",
   894 => x"64697265",
   895 => x"63746f72",
   896 => x"79207365",
   897 => x"63746f72",
   898 => x"2025640a",
   899 => x"00000000",
   900 => x"47657446",
   901 => x"41544c69",
   902 => x"6e6b2072",
   903 => x"65747572",
   904 => x"6e656420",
   905 => x"25640a00",
   906 => x"4f70656e",
   907 => x"65642066",
   908 => x"696c652c",
   909 => x"206c6f61",
   910 => x"64696e67",
   911 => x"2e2e2e0a",
   912 => x"00000000",
   913 => x"43616e27",
   914 => x"74206f70",
   915 => x"656e2025",
   916 => x"730a0000",
   917 => x"436d645f",
   918 => x"696e6974",
   919 => x"0a000000",
   920 => x"636d645f",
   921 => x"434d4438",
   922 => x"20726573",
   923 => x"706f6e73",
   924 => x"653a2025",
   925 => x"640a0000",
   926 => x"434d4438",
   927 => x"5f342072",
   928 => x"6573706f",
   929 => x"6e73653a",
   930 => x"2025640a",
   931 => x"00000000",
   932 => x"53444843",
   933 => x"20496e69",
   934 => x"7469616c",
   935 => x"697a6174",
   936 => x"696f6e20",
   937 => x"6572726f",
   938 => x"72210a00",
   939 => x"434d4435",
   940 => x"38202564",
   941 => x"0a202000",
   942 => x"434d4435",
   943 => x"385f3220",
   944 => x"25640a20",
   945 => x"20000000",
   946 => x"53504920",
   947 => x"496e6974",
   948 => x"28290a00",
   949 => x"52656164",
   950 => x"20636f6d",
   951 => x"6d616e64",
   952 => x"20666169",
   953 => x"6c656420",
   954 => x"61742025",
   955 => x"64202825",
   956 => x"64290a00",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

