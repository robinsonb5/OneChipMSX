-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b0bb1",
     9 => x"d0080b0b",
    10 => x"0bb1d408",
    11 => x"0b0b0bb1",
    12 => x"d8080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"b1d80c0b",
    16 => x"0b0bb1d4",
    17 => x"0c0b0b0b",
    18 => x"b1d00c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0ba8ac",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"b1d070b7",
    57 => x"ac278b38",
    58 => x"80717084",
    59 => x"05530c81",
    60 => x"e2048c51",
    61 => x"8aef0402",
    62 => x"fc050df8",
    63 => x"80518f0b",
    64 => x"b1e00c9f",
    65 => x"0bb1e40c",
    66 => x"a0717081",
    67 => x"055334b1",
    68 => x"e408ff05",
    69 => x"b1e40cb1",
    70 => x"e4088025",
    71 => x"eb38b1e0",
    72 => x"08ff05b1",
    73 => x"e00cb1e0",
    74 => x"088025d7",
    75 => x"38028405",
    76 => x"0d0402f0",
    77 => x"050df880",
    78 => x"53f8a054",
    79 => x"83bf5273",
    80 => x"70810555",
    81 => x"33517073",
    82 => x"70810555",
    83 => x"34ff1252",
    84 => x"718025eb",
    85 => x"38fbc053",
    86 => x"9f52a073",
    87 => x"70810555",
    88 => x"34ff1252",
    89 => x"718025f2",
    90 => x"38029005",
    91 => x"0d0402f4",
    92 => x"050d7453",
    93 => x"8e0bb1e0",
    94 => x"08258f38",
    95 => x"82b22db1",
    96 => x"e008ff05",
    97 => x"b1e00c82",
    98 => x"f404b1e0",
    99 => x"08b1e408",
   100 => x"5351728a",
   101 => x"2e098106",
   102 => x"b7387151",
   103 => x"719f24a0",
   104 => x"38b1e008",
   105 => x"a02911f8",
   106 => x"80115151",
   107 => x"a07134b1",
   108 => x"e4088105",
   109 => x"b1e40cb1",
   110 => x"e408519f",
   111 => x"7125e238",
   112 => x"800bb1e4",
   113 => x"0cb1e008",
   114 => x"8105b1e0",
   115 => x"0c83e404",
   116 => x"70a02912",
   117 => x"f8801151",
   118 => x"51727134",
   119 => x"b1e40881",
   120 => x"05b1e40c",
   121 => x"b1e408a0",
   122 => x"2e098106",
   123 => x"8e38800b",
   124 => x"b1e40cb1",
   125 => x"e0088105",
   126 => x"b1e00c02",
   127 => x"8c050d04",
   128 => x"02e8050d",
   129 => x"77795656",
   130 => x"880bfc16",
   131 => x"77712c8f",
   132 => x"06545254",
   133 => x"80537272",
   134 => x"25953871",
   135 => x"53fbe014",
   136 => x"51877134",
   137 => x"8114ff14",
   138 => x"545472f1",
   139 => x"387153f9",
   140 => x"1576712c",
   141 => x"87065351",
   142 => x"71802e8b",
   143 => x"38fbe014",
   144 => x"51717134",
   145 => x"81145472",
   146 => x"8e249538",
   147 => x"8f733153",
   148 => x"fbe01451",
   149 => x"a0713481",
   150 => x"14ff1454",
   151 => x"5472f138",
   152 => x"0298050d",
   153 => x"0402ec05",
   154 => x"0d800bb1",
   155 => x"e80cf68c",
   156 => x"08f69008",
   157 => x"71882c56",
   158 => x"5481ff06",
   159 => x"52737225",
   160 => x"88387154",
   161 => x"820bb1e8",
   162 => x"0c72882c",
   163 => x"7381ff06",
   164 => x"54557473",
   165 => x"258b3872",
   166 => x"b1e80884",
   167 => x"07b1e80c",
   168 => x"5573842b",
   169 => x"86a07125",
   170 => x"83713170",
   171 => x"0b0b0baf",
   172 => x"b40c8171",
   173 => x"2bff05f6",
   174 => x"880cfecc",
   175 => x"13ff122c",
   176 => x"788829ff",
   177 => x"94057081",
   178 => x"2cb1e808",
   179 => x"52585255",
   180 => x"51525476",
   181 => x"802e8538",
   182 => x"70810751",
   183 => x"70f6940c",
   184 => x"71098105",
   185 => x"f6800c72",
   186 => x"098105f6",
   187 => x"840c0294",
   188 => x"050d0402",
   189 => x"f4050d74",
   190 => x"53727081",
   191 => x"055480f5",
   192 => x"2d527180",
   193 => x"2e893871",
   194 => x"5182ee2d",
   195 => x"85f90402",
   196 => x"8c050d04",
   197 => x"02f8050d",
   198 => x"a2842d80",
   199 => x"da51a3bb",
   200 => x"2db1d008",
   201 => x"812a7081",
   202 => x"06515271",
   203 => x"802ee938",
   204 => x"0288050d",
   205 => x"0402f405",
   206 => x"0db79c08",
   207 => x"81c406b0",
   208 => x"b80b80f5",
   209 => x"2d525270",
   210 => x"802e8638",
   211 => x"71848007",
   212 => x"52aff00b",
   213 => x"80f52d72",
   214 => x"07b0880b",
   215 => x"80f52d70",
   216 => x"812a7081",
   217 => x"06515354",
   218 => x"5270802e",
   219 => x"86387182",
   220 => x"80075272",
   221 => x"81065170",
   222 => x"802e8538",
   223 => x"71880752",
   224 => x"b0940b80",
   225 => x"f52d7084",
   226 => x"2b730784",
   227 => x"32b1d00c",
   228 => x"51028c05",
   229 => x"0d0402f4",
   230 => x"050d7470",
   231 => x"8432b79c",
   232 => x"0c708306",
   233 => x"525370af",
   234 => x"e80b8805",
   235 => x"81b72d72",
   236 => x"892a7081",
   237 => x"06515170",
   238 => x"b0b80b81",
   239 => x"b72d7283",
   240 => x"2a810673",
   241 => x"882a7081",
   242 => x"06515252",
   243 => x"70802e85",
   244 => x"38718207",
   245 => x"5271b088",
   246 => x"0b81b72d",
   247 => x"72842c70",
   248 => x"83065151",
   249 => x"70b0940b",
   250 => x"81b72d70",
   251 => x"b1d00c02",
   252 => x"8c050d04",
   253 => x"02d4050d",
   254 => x"aaf85185",
   255 => x"f32d9a85",
   256 => x"2db1d008",
   257 => x"802e82ab",
   258 => x"3886b52d",
   259 => x"b1d00853",
   260 => x"8ce02db1",
   261 => x"d00854b1",
   262 => x"d008802e",
   263 => x"8297389c",
   264 => x"c82db1d0",
   265 => x"08802e87",
   266 => x"38ab9051",
   267 => x"88bc0495",
   268 => x"e72db1d0",
   269 => x"08802e9c",
   270 => x"38abd051",
   271 => x"85f32d86",
   272 => x"942d7284",
   273 => x"0753810b",
   274 => x"fec40c72",
   275 => x"fec00c72",
   276 => x"5187962d",
   277 => x"840bfec4",
   278 => x"0cac9851",
   279 => x"85f32dac",
   280 => x"b052b1f0",
   281 => x"5192fc2d",
   282 => x"b1d00898",
   283 => x"38acbc51",
   284 => x"85f32dac",
   285 => x"d452b1f0",
   286 => x"5192fc2d",
   287 => x"b1d00880",
   288 => x"2e81b038",
   289 => x"ace05185",
   290 => x"f32db1f4",
   291 => x"08578077",
   292 => x"595a767a",
   293 => x"2e8b3881",
   294 => x"1a78812a",
   295 => x"595a77f7",
   296 => x"38f71a5a",
   297 => x"80772581",
   298 => x"80387952",
   299 => x"77518480",
   300 => x"2db1fc52",
   301 => x"b1f05195",
   302 => x"c12db1d0",
   303 => x"0853b1d0",
   304 => x"08802e80",
   305 => x"c938b1fc",
   306 => x"5b805989",
   307 => x"fb047a70",
   308 => x"84055c08",
   309 => x"7081ff06",
   310 => x"71882c70",
   311 => x"81ff0673",
   312 => x"902c7081",
   313 => x"ff067598",
   314 => x"2afec80c",
   315 => x"fec80c58",
   316 => x"fec80c57",
   317 => x"fec80c84",
   318 => x"1a5a5376",
   319 => x"53848077",
   320 => x"25843884",
   321 => x"80537279",
   322 => x"24c4388a",
   323 => x"9904acfc",
   324 => x"5185f32d",
   325 => x"72548ab5",
   326 => x"04b1f051",
   327 => x"95942dfc",
   328 => x"80178119",
   329 => x"595789a4",
   330 => x"04820bfe",
   331 => x"c40c8154",
   332 => x"8ab50480",
   333 => x"5473b1d0",
   334 => x"0c02ac05",
   335 => x"0d0402f8",
   336 => x"050da48b",
   337 => x"2d81f72d",
   338 => x"815184e5",
   339 => x"2dfec452",
   340 => x"81720ca1",
   341 => x"d12da1d1",
   342 => x"2d84720c",
   343 => x"87f42daf",
   344 => x"b851a5a4",
   345 => x"2d805184",
   346 => x"e52d0288",
   347 => x"050d0402",
   348 => x"f4050d84",
   349 => x"b9518796",
   350 => x"2d810bfe",
   351 => x"c40c84b9",
   352 => x"0bfec00c",
   353 => x"840bfec4",
   354 => x"0ca1ec2d",
   355 => x"a3ff2da1",
   356 => x"d12da1d1",
   357 => x"2d81f72d",
   358 => x"815184e5",
   359 => x"2da1d12d",
   360 => x"a1d12d81",
   361 => x"5184e52d",
   362 => x"87f42db1",
   363 => x"d008802e",
   364 => x"80db3880",
   365 => x"5184e52d",
   366 => x"afb851a5",
   367 => x"a42da284",
   368 => x"2da5b42d",
   369 => x"b1d00853",
   370 => x"86b52db1",
   371 => x"d008fec0",
   372 => x"0c86b52d",
   373 => x"b1d008b1",
   374 => x"ec082e9c",
   375 => x"38b1d008",
   376 => x"b1ec0c85",
   377 => x"52725184",
   378 => x"e52da1d1",
   379 => x"2da1d12d",
   380 => x"ff125271",
   381 => x"8025ee38",
   382 => x"72802e89",
   383 => x"388a0bfe",
   384 => x"c40c8bbe",
   385 => x"04820bfe",
   386 => x"c40c8bbe",
   387 => x"04ad9051",
   388 => x"85f32d82",
   389 => x"0bfec40c",
   390 => x"800bb1d0",
   391 => x"0c028c05",
   392 => x"0d0402e8",
   393 => x"050d7779",
   394 => x"7b585555",
   395 => x"80537276",
   396 => x"25a33874",
   397 => x"70810556",
   398 => x"80f52d74",
   399 => x"70810556",
   400 => x"80f52d52",
   401 => x"5271712e",
   402 => x"86388151",
   403 => x"8cd70481",
   404 => x"13538cae",
   405 => x"04805170",
   406 => x"b1d00c02",
   407 => x"98050d04",
   408 => x"02d8050d",
   409 => x"800bb684",
   410 => x"0cb1fc52",
   411 => x"80519ba5",
   412 => x"2db1d008",
   413 => x"54b1d008",
   414 => x"8c38ada8",
   415 => x"5185f32d",
   416 => x"73559285",
   417 => x"04805681",
   418 => x"0bb6a80c",
   419 => x"8853adbc",
   420 => x"52b2b251",
   421 => x"8ca22db1",
   422 => x"d008762e",
   423 => x"09810687",
   424 => x"38b1d008",
   425 => x"b6a80c88",
   426 => x"53adc852",
   427 => x"b2ce518c",
   428 => x"a22db1d0",
   429 => x"088738b1",
   430 => x"d008b6a8",
   431 => x"0cb6a808",
   432 => x"52add451",
   433 => x"9ec22db6",
   434 => x"a808802e",
   435 => x"80f638b5",
   436 => x"c20b80f5",
   437 => x"2db5c30b",
   438 => x"80f52d71",
   439 => x"982b7190",
   440 => x"2b07b5c4",
   441 => x"0b80f52d",
   442 => x"70882b72",
   443 => x"07b5c50b",
   444 => x"80f52d71",
   445 => x"07b5fa0b",
   446 => x"80f52db5",
   447 => x"fb0b80f5",
   448 => x"2d71882b",
   449 => x"07535f54",
   450 => x"525a5657",
   451 => x"557381ab",
   452 => x"aa2e0981",
   453 => x"068d3875",
   454 => x"519d972d",
   455 => x"b1d00856",
   456 => x"8eb00473",
   457 => x"82d4d52e",
   458 => x"8738adec",
   459 => x"518ef104",
   460 => x"b1fc5275",
   461 => x"519ba52d",
   462 => x"b1d00855",
   463 => x"b1d00880",
   464 => x"2e83c238",
   465 => x"8853adc8",
   466 => x"52b2ce51",
   467 => x"8ca22db1",
   468 => x"d0088938",
   469 => x"810bb684",
   470 => x"0c8ef704",
   471 => x"8853adbc",
   472 => x"52b2b251",
   473 => x"8ca22db1",
   474 => x"d008802e",
   475 => x"8a38ae8c",
   476 => x"5185f32d",
   477 => x"8fd104b5",
   478 => x"fa0b80f5",
   479 => x"2d547380",
   480 => x"d52e0981",
   481 => x"0680ca38",
   482 => x"b5fb0b80",
   483 => x"f52d5473",
   484 => x"81aa2e09",
   485 => x"8106ba38",
   486 => x"800bb1fc",
   487 => x"0b80f52d",
   488 => x"56547481",
   489 => x"e92e8338",
   490 => x"81547481",
   491 => x"eb2e8c38",
   492 => x"80557375",
   493 => x"2e098106",
   494 => x"82cb38b2",
   495 => x"870b80f5",
   496 => x"2d55748d",
   497 => x"38b2880b",
   498 => x"80f52d54",
   499 => x"73822e86",
   500 => x"38805592",
   501 => x"8504b289",
   502 => x"0b80f52d",
   503 => x"70b5fc0c",
   504 => x"ff05b680",
   505 => x"0cb28a0b",
   506 => x"80f52db2",
   507 => x"8b0b80f5",
   508 => x"2d587605",
   509 => x"77828029",
   510 => x"0570b688",
   511 => x"0cb28c0b",
   512 => x"80f52d70",
   513 => x"b69c0cb6",
   514 => x"84085957",
   515 => x"5876802e",
   516 => x"81a33888",
   517 => x"53adc852",
   518 => x"b2ce518c",
   519 => x"a22db1d0",
   520 => x"0881e238",
   521 => x"b5fc0870",
   522 => x"842bb6a0",
   523 => x"0c70b698",
   524 => x"0cb2a10b",
   525 => x"80f52db2",
   526 => x"a00b80f5",
   527 => x"2d718280",
   528 => x"2905b2a2",
   529 => x"0b80f52d",
   530 => x"70848080",
   531 => x"2912b2a3",
   532 => x"0b80f52d",
   533 => x"7081800a",
   534 => x"291270b6",
   535 => x"a40cb69c",
   536 => x"087129b6",
   537 => x"88080570",
   538 => x"b68c0cb2",
   539 => x"a90b80f5",
   540 => x"2db2a80b",
   541 => x"80f52d71",
   542 => x"82802905",
   543 => x"b2aa0b80",
   544 => x"f52d7084",
   545 => x"80802912",
   546 => x"b2ab0b80",
   547 => x"f52d7098",
   548 => x"2b81f00a",
   549 => x"06720570",
   550 => x"b6900cfe",
   551 => x"117e2977",
   552 => x"05b6940c",
   553 => x"52595243",
   554 => x"545e5152",
   555 => x"59525d57",
   556 => x"59579283",
   557 => x"04b28e0b",
   558 => x"80f52db2",
   559 => x"8d0b80f5",
   560 => x"2d718280",
   561 => x"290570b6",
   562 => x"a00c70a0",
   563 => x"2983ff05",
   564 => x"70892a70",
   565 => x"b6980cb2",
   566 => x"930b80f5",
   567 => x"2db2920b",
   568 => x"80f52d71",
   569 => x"82802905",
   570 => x"70b6a40c",
   571 => x"7b71291e",
   572 => x"70b6940c",
   573 => x"7db6900c",
   574 => x"7305b68c",
   575 => x"0c555e51",
   576 => x"51555581",
   577 => x"5574b1d0",
   578 => x"0c02a805",
   579 => x"0d0402ec",
   580 => x"050d7670",
   581 => x"872c7180",
   582 => x"ff065556",
   583 => x"54b68408",
   584 => x"8a387388",
   585 => x"2c7481ff",
   586 => x"065455b1",
   587 => x"fc52b688",
   588 => x"0815519b",
   589 => x"a52db1d0",
   590 => x"0854b1d0",
   591 => x"08802eb3",
   592 => x"38b68408",
   593 => x"802e9838",
   594 => x"728429b1",
   595 => x"fc057008",
   596 => x"52539d97",
   597 => x"2db1d008",
   598 => x"f00a0653",
   599 => x"92f10472",
   600 => x"10b1fc05",
   601 => x"7080e02d",
   602 => x"52539dc7",
   603 => x"2db1d008",
   604 => x"53725473",
   605 => x"b1d00c02",
   606 => x"94050d04",
   607 => x"02c8050d",
   608 => x"7f615f5b",
   609 => x"800bb690",
   610 => x"08b69408",
   611 => x"595d56b6",
   612 => x"8408762e",
   613 => x"8a38b5fc",
   614 => x"08842b58",
   615 => x"93a504b6",
   616 => x"9808842b",
   617 => x"58805978",
   618 => x"782781a9",
   619 => x"38788f06",
   620 => x"a0175754",
   621 => x"738f38b1",
   622 => x"fc527651",
   623 => x"8117579b",
   624 => x"a52db1fc",
   625 => x"56807680",
   626 => x"f52d5654",
   627 => x"74742e83",
   628 => x"38815474",
   629 => x"81e52e80",
   630 => x"f6388170",
   631 => x"7506555d",
   632 => x"73802e80",
   633 => x"ea388b16",
   634 => x"80f52d98",
   635 => x"065a7980",
   636 => x"de388b53",
   637 => x"7d527551",
   638 => x"8ca22db1",
   639 => x"d00880cf",
   640 => x"389c1608",
   641 => x"519d972d",
   642 => x"b1d00884",
   643 => x"1c0c9a16",
   644 => x"80e02d51",
   645 => x"9dc72db1",
   646 => x"d008b1d0",
   647 => x"08881d0c",
   648 => x"b1d00855",
   649 => x"55b68408",
   650 => x"802e9838",
   651 => x"941680e0",
   652 => x"2d519dc7",
   653 => x"2db1d008",
   654 => x"902b83ff",
   655 => x"f00a0670",
   656 => x"16515473",
   657 => x"881c0c79",
   658 => x"7b0c7c54",
   659 => x"958b0481",
   660 => x"195993a7",
   661 => x"04b68408",
   662 => x"802eae38",
   663 => x"7b51928e",
   664 => x"2db1d008",
   665 => x"b1d00880",
   666 => x"fffffff8",
   667 => x"06555c73",
   668 => x"80ffffff",
   669 => x"f82e9238",
   670 => x"b1d008fe",
   671 => x"05b5fc08",
   672 => x"29b68c08",
   673 => x"055793a5",
   674 => x"04805473",
   675 => x"b1d00c02",
   676 => x"b8050d04",
   677 => x"02f4050d",
   678 => x"74700881",
   679 => x"05710c70",
   680 => x"08b68008",
   681 => x"06535371",
   682 => x"8e388813",
   683 => x"0851928e",
   684 => x"2db1d008",
   685 => x"88140c81",
   686 => x"0bb1d00c",
   687 => x"028c050d",
   688 => x"0402f005",
   689 => x"0d758811",
   690 => x"08fe05b5",
   691 => x"fc0829b6",
   692 => x"8c081172",
   693 => x"08b68008",
   694 => x"06057955",
   695 => x"5354549b",
   696 => x"a52d0290",
   697 => x"050d04b6",
   698 => x"8408b1d0",
   699 => x"0c0402f4",
   700 => x"050dd452",
   701 => x"81ff720c",
   702 => x"71085381",
   703 => x"ff720c72",
   704 => x"882b83fe",
   705 => x"80067208",
   706 => x"7081ff06",
   707 => x"51525381",
   708 => x"ff720c72",
   709 => x"7107882b",
   710 => x"72087081",
   711 => x"ff065152",
   712 => x"5381ff72",
   713 => x"0c727107",
   714 => x"882b7208",
   715 => x"7081ff06",
   716 => x"7207b1d0",
   717 => x"0c525302",
   718 => x"8c050d04",
   719 => x"02f4050d",
   720 => x"74767181",
   721 => x"ff06d40c",
   722 => x"5353b6ac",
   723 => x"08853871",
   724 => x"892b5271",
   725 => x"982ad40c",
   726 => x"71902a70",
   727 => x"81ff06d4",
   728 => x"0c517188",
   729 => x"2a7081ff",
   730 => x"06d40c51",
   731 => x"7181ff06",
   732 => x"d40c7290",
   733 => x"2a7081ff",
   734 => x"06d40c51",
   735 => x"d4087081",
   736 => x"ff065151",
   737 => x"82b8bf52",
   738 => x"7081ff2e",
   739 => x"09810694",
   740 => x"3881ff0b",
   741 => x"d40cd408",
   742 => x"7081ff06",
   743 => x"ff145451",
   744 => x"5171e538",
   745 => x"70b1d00c",
   746 => x"028c050d",
   747 => x"0402fc05",
   748 => x"0d81c751",
   749 => x"81ff0bd4",
   750 => x"0cff1151",
   751 => x"708025f4",
   752 => x"38028405",
   753 => x"0d0402f0",
   754 => x"050d97ad",
   755 => x"2d8fcf53",
   756 => x"805287fc",
   757 => x"80f75196",
   758 => x"bc2db1d0",
   759 => x"0854b1d0",
   760 => x"08812e09",
   761 => x"8106a338",
   762 => x"81ff0bd4",
   763 => x"0c820a52",
   764 => x"849c80e9",
   765 => x"5196bc2d",
   766 => x"b1d0088b",
   767 => x"3881ff0b",
   768 => x"d40c7353",
   769 => x"98900497",
   770 => x"ad2dff13",
   771 => x"5372c138",
   772 => x"72b1d00c",
   773 => x"0290050d",
   774 => x"0402f405",
   775 => x"0d81ff0b",
   776 => x"d40c9353",
   777 => x"805287fc",
   778 => x"80c15196",
   779 => x"bc2db1d0",
   780 => x"088b3881",
   781 => x"ff0bd40c",
   782 => x"815398c6",
   783 => x"0497ad2d",
   784 => x"ff135372",
   785 => x"df3872b1",
   786 => x"d00c028c",
   787 => x"050d0402",
   788 => x"f0050d97",
   789 => x"ad2d83aa",
   790 => x"52849c80",
   791 => x"c85196bc",
   792 => x"2db1d008",
   793 => x"812e0981",
   794 => x"06923895",
   795 => x"ee2db1d0",
   796 => x"0883ffff",
   797 => x"06537283",
   798 => x"aa2e9738",
   799 => x"98992d99",
   800 => x"8d048154",
   801 => x"99fc04ae",
   802 => x"ac5185f3",
   803 => x"2d805499",
   804 => x"fc0481ff",
   805 => x"0bd40cb1",
   806 => x"5397c62d",
   807 => x"b1d00880",
   808 => x"2e80ca38",
   809 => x"805287fc",
   810 => x"80fa5196",
   811 => x"bc2db1d0",
   812 => x"08b13881",
   813 => x"ff0bd40c",
   814 => x"d4085381",
   815 => x"ff0bd40c",
   816 => x"81ff0bd4",
   817 => x"0c81ff0b",
   818 => x"d40c81ff",
   819 => x"0bd40c72",
   820 => x"862a7081",
   821 => x"06b1d008",
   822 => x"56515372",
   823 => x"802e9d38",
   824 => x"998204b1",
   825 => x"d00852ae",
   826 => x"c8519ec2",
   827 => x"2d72822e",
   828 => x"ff9538ff",
   829 => x"135372ff",
   830 => x"a0387254",
   831 => x"73b1d00c",
   832 => x"0290050d",
   833 => x"0402f405",
   834 => x"0d810bb6",
   835 => x"ac0cd008",
   836 => x"708f2a70",
   837 => x"81065151",
   838 => x"5372f338",
   839 => x"72d00c97",
   840 => x"ad2daed4",
   841 => x"5185f32d",
   842 => x"d008708f",
   843 => x"2a708106",
   844 => x"51515372",
   845 => x"f338810b",
   846 => x"d00c80e3",
   847 => x"53805284",
   848 => x"d480c051",
   849 => x"96bc2db1",
   850 => x"d008812e",
   851 => x"9a387282",
   852 => x"2e098106",
   853 => x"8c38aef0",
   854 => x"5185f32d",
   855 => x"80539b9c",
   856 => x"04ff1353",
   857 => x"72d73898",
   858 => x"cf2db1d0",
   859 => x"08b6ac0c",
   860 => x"b1d0088b",
   861 => x"38815287",
   862 => x"fc80d051",
   863 => x"96bc2d81",
   864 => x"ff0bd40c",
   865 => x"d008708f",
   866 => x"2a708106",
   867 => x"51515372",
   868 => x"f33872d0",
   869 => x"0c81ff0b",
   870 => x"d40c8153",
   871 => x"72b1d00c",
   872 => x"028c050d",
   873 => x"0402e005",
   874 => x"0d797b57",
   875 => x"57805881",
   876 => x"ff0bd40c",
   877 => x"d008708f",
   878 => x"2a708106",
   879 => x"51515473",
   880 => x"f3388281",
   881 => x"0bd00c81",
   882 => x"ff0bd40c",
   883 => x"765287fc",
   884 => x"80d15196",
   885 => x"bc2d80db",
   886 => x"c6df55b1",
   887 => x"d008802e",
   888 => x"9038b1d0",
   889 => x"08537652",
   890 => x"af88519e",
   891 => x"c22d9cbf",
   892 => x"0481ff0b",
   893 => x"d40cd408",
   894 => x"7081ff06",
   895 => x"51547381",
   896 => x"fe2e0981",
   897 => x"069d3880",
   898 => x"ff5495ee",
   899 => x"2db1d008",
   900 => x"76708405",
   901 => x"580cff14",
   902 => x"54738025",
   903 => x"ed388158",
   904 => x"9ca904ff",
   905 => x"155574c9",
   906 => x"3881ff0b",
   907 => x"d40cd008",
   908 => x"708f2a70",
   909 => x"81065151",
   910 => x"5473f338",
   911 => x"73d00c77",
   912 => x"b1d00c02",
   913 => x"a0050d04",
   914 => x"b6ac08b1",
   915 => x"d00c0402",
   916 => x"e8050d80",
   917 => x"78575575",
   918 => x"70840557",
   919 => x"08538054",
   920 => x"72982a73",
   921 => x"882b5452",
   922 => x"71802ea2",
   923 => x"38c00870",
   924 => x"882a7081",
   925 => x"06515151",
   926 => x"70802ef1",
   927 => x"3871c00c",
   928 => x"81158115",
   929 => x"55558374",
   930 => x"25d63871",
   931 => x"ca3874b1",
   932 => x"d00c0298",
   933 => x"050d0402",
   934 => x"f4050d74",
   935 => x"70882a83",
   936 => x"fe800670",
   937 => x"72982a07",
   938 => x"72882b87",
   939 => x"fc808006",
   940 => x"73982b81",
   941 => x"f00a0671",
   942 => x"730707b1",
   943 => x"d00c5651",
   944 => x"5351028c",
   945 => x"050d0402",
   946 => x"f8050d02",
   947 => x"8e0580f5",
   948 => x"2d74882b",
   949 => x"077083ff",
   950 => x"ff06b1d0",
   951 => x"0c510288",
   952 => x"050d0402",
   953 => x"ec050d76",
   954 => x"53805572",
   955 => x"75258b38",
   956 => x"ad5182ee",
   957 => x"2d720981",
   958 => x"05537280",
   959 => x"2eb53887",
   960 => x"54729c2a",
   961 => x"73842b54",
   962 => x"5271802e",
   963 => x"83388155",
   964 => x"89722587",
   965 => x"38b71252",
   966 => x"9e9e04b0",
   967 => x"12527480",
   968 => x"2e863871",
   969 => x"5182ee2d",
   970 => x"ff145473",
   971 => x"8025d238",
   972 => x"9eb804b0",
   973 => x"5182ee2d",
   974 => x"800bb1d0",
   975 => x"0c029405",
   976 => x"0d0402c0",
   977 => x"050d0280",
   978 => x"c4055780",
   979 => x"70787084",
   980 => x"055a0872",
   981 => x"415f5d58",
   982 => x"7c708405",
   983 => x"5e085a80",
   984 => x"5b79982a",
   985 => x"7a882b5b",
   986 => x"56758638",
   987 => x"775fa0ba",
   988 => x"047d802e",
   989 => x"81a23880",
   990 => x"5e7580e4",
   991 => x"2e8a3875",
   992 => x"80f82e09",
   993 => x"81068938",
   994 => x"76841871",
   995 => x"085e5854",
   996 => x"7580e42e",
   997 => x"9f387580",
   998 => x"e4268a38",
   999 => x"7580e32e",
  1000 => x"be389fea",
  1001 => x"047580f3",
  1002 => x"2ea33875",
  1003 => x"80f82e89",
  1004 => x"389fea04",
  1005 => x"8a539fbb",
  1006 => x"049053b6",
  1007 => x"b0527b51",
  1008 => x"9de32db1",
  1009 => x"d008b6b0",
  1010 => x"5a559ffa",
  1011 => x"04768418",
  1012 => x"71087054",
  1013 => x"5b58549c",
  1014 => x"cf2d8055",
  1015 => x"9ffa0476",
  1016 => x"84187108",
  1017 => x"585854a0",
  1018 => x"a504a551",
  1019 => x"82ee2d75",
  1020 => x"5182ee2d",
  1021 => x"821858a0",
  1022 => x"ad0474ff",
  1023 => x"16565480",
  1024 => x"7425aa38",
  1025 => x"78708105",
  1026 => x"5a80f52d",
  1027 => x"70525682",
  1028 => x"ee2d8118",
  1029 => x"589ffa04",
  1030 => x"75a52e09",
  1031 => x"81068638",
  1032 => x"815ea0ad",
  1033 => x"04755182",
  1034 => x"ee2d8118",
  1035 => x"58811b5b",
  1036 => x"837b25fe",
  1037 => x"ac3875fe",
  1038 => x"9f387eb1",
  1039 => x"d00c0280",
  1040 => x"c0050d04",
  1041 => x"02fc050d",
  1042 => x"72518071",
  1043 => x"0c800b84",
  1044 => x"120c0284",
  1045 => x"050d0402",
  1046 => x"f0050d75",
  1047 => x"70088412",
  1048 => x"08535353",
  1049 => x"ff547171",
  1050 => x"2e9b3884",
  1051 => x"13087084",
  1052 => x"29148b11",
  1053 => x"80f52d84",
  1054 => x"16088111",
  1055 => x"87068418",
  1056 => x"0c525651",
  1057 => x"5173b1d0",
  1058 => x"0c029005",
  1059 => x"0d0402f8",
  1060 => x"050da485",
  1061 => x"2de00870",
  1062 => x"8b2a7081",
  1063 => x"06515252",
  1064 => x"70802e9d",
  1065 => x"38b6f008",
  1066 => x"708429b6",
  1067 => x"f8057381",
  1068 => x"ff06710c",
  1069 => x"5151b6f0",
  1070 => x"08811187",
  1071 => x"06b6f00c",
  1072 => x"51800bb7",
  1073 => x"980ca3f8",
  1074 => x"2da3ff2d",
  1075 => x"0288050d",
  1076 => x"0402fc05",
  1077 => x"0da4852d",
  1078 => x"810bb798",
  1079 => x"0ca3ff2d",
  1080 => x"b7980851",
  1081 => x"70fa3802",
  1082 => x"84050d04",
  1083 => x"02fc050d",
  1084 => x"b6f051a0",
  1085 => x"c42da18e",
  1086 => x"51a3f42d",
  1087 => x"a39e2d02",
  1088 => x"84050d04",
  1089 => x"02f4050d",
  1090 => x"a38604b1",
  1091 => x"d00881f0",
  1092 => x"2e098106",
  1093 => x"8938810b",
  1094 => x"b1c40ca3",
  1095 => x"8604b1d0",
  1096 => x"0881e02e",
  1097 => x"09810689",
  1098 => x"38810bb1",
  1099 => x"c80ca386",
  1100 => x"04b1d008",
  1101 => x"52b1c808",
  1102 => x"802e8838",
  1103 => x"b1d00881",
  1104 => x"80055271",
  1105 => x"842c728f",
  1106 => x"065353b1",
  1107 => x"c408802e",
  1108 => x"99387284",
  1109 => x"29b18405",
  1110 => x"72138171",
  1111 => x"2b700973",
  1112 => x"0806730c",
  1113 => x"515353a2",
  1114 => x"fc047284",
  1115 => x"29b18405",
  1116 => x"72138371",
  1117 => x"2b720807",
  1118 => x"720c5353",
  1119 => x"800bb1c8",
  1120 => x"0c800bb1",
  1121 => x"c40cb6f0",
  1122 => x"51a0d72d",
  1123 => x"b1d008ff",
  1124 => x"24fef838",
  1125 => x"800bb1d0",
  1126 => x"0c028c05",
  1127 => x"0d0402f8",
  1128 => x"050db184",
  1129 => x"528f5180",
  1130 => x"72708405",
  1131 => x"540cff11",
  1132 => x"51708025",
  1133 => x"f2380288",
  1134 => x"050d0402",
  1135 => x"f0050d75",
  1136 => x"51a4852d",
  1137 => x"70822cfc",
  1138 => x"06b18411",
  1139 => x"72109e06",
  1140 => x"71087072",
  1141 => x"2a708306",
  1142 => x"82742b70",
  1143 => x"09740676",
  1144 => x"0c545156",
  1145 => x"57535153",
  1146 => x"a3ff2d71",
  1147 => x"b1d00c02",
  1148 => x"90050d04",
  1149 => x"71980c04",
  1150 => x"ffb008b1",
  1151 => x"d00c0481",
  1152 => x"0bffb00c",
  1153 => x"04800bff",
  1154 => x"b00c0402",
  1155 => x"fc050d80",
  1156 => x"0bb1cc0c",
  1157 => x"805184e5",
  1158 => x"2d028405",
  1159 => x"0d0402f0",
  1160 => x"050db7a0",
  1161 => x"085481f7",
  1162 => x"2d800bb7",
  1163 => x"a40c7308",
  1164 => x"802e80eb",
  1165 => x"38820bb1",
  1166 => x"e40cb7a4",
  1167 => x"088f06b1",
  1168 => x"e00c7308",
  1169 => x"5271812e",
  1170 => x"a4387183",
  1171 => x"2e098106",
  1172 => x"b9388814",
  1173 => x"80f52d84",
  1174 => x"1508afa8",
  1175 => x"53545285",
  1176 => x"f32d7184",
  1177 => x"29137008",
  1178 => x"5252a58e",
  1179 => x"04b79c08",
  1180 => x"8815082c",
  1181 => x"70810651",
  1182 => x"5271802e",
  1183 => x"8738afac",
  1184 => x"51a58704",
  1185 => x"afb05185",
  1186 => x"f32d8414",
  1187 => x"085185f3",
  1188 => x"2db7a408",
  1189 => x"8105b7a4",
  1190 => x"0c8c1454",
  1191 => x"a4ae0402",
  1192 => x"90050d04",
  1193 => x"71b7a00c",
  1194 => x"a49e2db7",
  1195 => x"a408ff05",
  1196 => x"b7a80c04",
  1197 => x"02f0050d",
  1198 => x"8751a3bb",
  1199 => x"2db1d008",
  1200 => x"812a7081",
  1201 => x"06515271",
  1202 => x"802ea038",
  1203 => x"a5d204a2",
  1204 => x"842d8751",
  1205 => x"a3bb2db1",
  1206 => x"d008f438",
  1207 => x"b1cc0881",
  1208 => x"3270b1cc",
  1209 => x"0c705252",
  1210 => x"84e52db1",
  1211 => x"cc089638",
  1212 => x"80da51a3",
  1213 => x"bb2d81f5",
  1214 => x"51a3bb2d",
  1215 => x"81f251a3",
  1216 => x"bb2da8a2",
  1217 => x"0481f551",
  1218 => x"a3bb2db1",
  1219 => x"d008812a",
  1220 => x"70810651",
  1221 => x"5271802e",
  1222 => x"8f38b7a8",
  1223 => x"08527180",
  1224 => x"2e8638ff",
  1225 => x"12b7a80c",
  1226 => x"81f251a3",
  1227 => x"bb2db1d0",
  1228 => x"08812a70",
  1229 => x"81065152",
  1230 => x"71802e95",
  1231 => x"38b7a408",
  1232 => x"ff05b7a8",
  1233 => x"08545272",
  1234 => x"72258638",
  1235 => x"8113b7a8",
  1236 => x"0c80da51",
  1237 => x"a3bb2db1",
  1238 => x"d008812a",
  1239 => x"70810651",
  1240 => x"5271802e",
  1241 => x"80fb38b7",
  1242 => x"a008b7a8",
  1243 => x"08555373",
  1244 => x"802e8a38",
  1245 => x"8c13ff15",
  1246 => x"5553a6ef",
  1247 => x"04720852",
  1248 => x"71822ea6",
  1249 => x"38718226",
  1250 => x"89387181",
  1251 => x"2ea538a7",
  1252 => x"e1047183",
  1253 => x"2ead3871",
  1254 => x"842e0981",
  1255 => x"0680c238",
  1256 => x"88130851",
  1257 => x"a5a42da7",
  1258 => x"e1048813",
  1259 => x"0852712d",
  1260 => x"a7e10481",
  1261 => x"0b881408",
  1262 => x"2bb79c08",
  1263 => x"32b79c0c",
  1264 => x"a7de0488",
  1265 => x"1380f52d",
  1266 => x"81058b14",
  1267 => x"80f52d53",
  1268 => x"54717424",
  1269 => x"83388054",
  1270 => x"73881481",
  1271 => x"b72da49e",
  1272 => x"2d805480",
  1273 => x"0bb1e40c",
  1274 => x"738f06b1",
  1275 => x"e00ca052",
  1276 => x"73b7a808",
  1277 => x"2e098106",
  1278 => x"9838b7a4",
  1279 => x"08ff0574",
  1280 => x"32700981",
  1281 => x"05707207",
  1282 => x"9f2a9171",
  1283 => x"31515153",
  1284 => x"53715182",
  1285 => x"ee2d8114",
  1286 => x"548e7425",
  1287 => x"c638b1cc",
  1288 => x"085271b1",
  1289 => x"d00c0290",
  1290 => x"050d0400",
  1291 => x"00ffffff",
  1292 => x"ff00ffff",
  1293 => x"ffff00ff",
  1294 => x"ffffff00",
  1295 => x"44495020",
  1296 => x"53776974",
  1297 => x"63686573",
  1298 => x"20100000",
  1299 => x"52657365",
  1300 => x"74000000",
  1301 => x"45786974",
  1302 => x"00000000",
  1303 => x"53442043",
  1304 => x"61726400",
  1305 => x"4a617061",
  1306 => x"6e657365",
  1307 => x"206b6579",
  1308 => x"626f6172",
  1309 => x"64206c61",
  1310 => x"796f7574",
  1311 => x"00000000",
  1312 => x"54757262",
  1313 => x"6f202831",
  1314 => x"302e3734",
  1315 => x"4d487a29",
  1316 => x"00000000",
  1317 => x"4261636b",
  1318 => x"00000000",
  1319 => x"32303438",
  1320 => x"4c422052",
  1321 => x"414d0000",
  1322 => x"34303936",
  1323 => x"4b422052",
  1324 => x"414d0000",
  1325 => x"536c323a",
  1326 => x"204e6f6e",
  1327 => x"65000000",
  1328 => x"536c323a",
  1329 => x"20455345",
  1330 => x"2d534343",
  1331 => x"20314d42",
  1332 => x"2f534343",
  1333 => x"2d490000",
  1334 => x"536c323a",
  1335 => x"20455345",
  1336 => x"2d52414d",
  1337 => x"20314d42",
  1338 => x"2f415343",
  1339 => x"49493800",
  1340 => x"536c323a",
  1341 => x"20455345",
  1342 => x"2d52414d",
  1343 => x"20314d42",
  1344 => x"2f415343",
  1345 => x"49493136",
  1346 => x"00000000",
  1347 => x"536c313a",
  1348 => x"204e6f6e",
  1349 => x"65000000",
  1350 => x"536c313a",
  1351 => x"20455345",
  1352 => x"2d534343",
  1353 => x"20314d42",
  1354 => x"2f534343",
  1355 => x"2d490000",
  1356 => x"536c313a",
  1357 => x"204d6567",
  1358 => x"6152414d",
  1359 => x"00000000",
  1360 => x"56474120",
  1361 => x"2d203331",
  1362 => x"4b487a2c",
  1363 => x"20363048",
  1364 => x"7a000000",
  1365 => x"56474120",
  1366 => x"2d203331",
  1367 => x"4b487a2c",
  1368 => x"20353048",
  1369 => x"7a000000",
  1370 => x"5456202d",
  1371 => x"20343830",
  1372 => x"692c2036",
  1373 => x"30487a00",
  1374 => x"496e6974",
  1375 => x"69616c69",
  1376 => x"7a696e67",
  1377 => x"20534420",
  1378 => x"63617264",
  1379 => x"0a000000",
  1380 => x"53444843",
  1381 => x"20636172",
  1382 => x"64206465",
  1383 => x"74656374",
  1384 => x"65642062",
  1385 => x"7574206e",
  1386 => x"6f740a73",
  1387 => x"7570706f",
  1388 => x"72746564",
  1389 => x"3b206469",
  1390 => x"7361626c",
  1391 => x"696e6720",
  1392 => x"53442063",
  1393 => x"6172640a",
  1394 => x"10204f4b",
  1395 => x"0a000000",
  1396 => x"46617433",
  1397 => x"32206669",
  1398 => x"6c657379",
  1399 => x"7374656d",
  1400 => x"20646574",
  1401 => x"65637465",
  1402 => x"64206275",
  1403 => x"740a6e6f",
  1404 => x"74207375",
  1405 => x"70706f72",
  1406 => x"7465643b",
  1407 => x"20646973",
  1408 => x"61626c69",
  1409 => x"6e672053",
  1410 => x"44206361",
  1411 => x"72640a10",
  1412 => x"204f4b0a",
  1413 => x"00000000",
  1414 => x"54727969",
  1415 => x"6e67204d",
  1416 => x"53583342",
  1417 => x"494f532e",
  1418 => x"5359532e",
  1419 => x"2e2e0a00",
  1420 => x"4d535833",
  1421 => x"42494f53",
  1422 => x"53595300",
  1423 => x"54727969",
  1424 => x"6e672042",
  1425 => x"494f535f",
  1426 => x"4d32502e",
  1427 => x"524f4d2e",
  1428 => x"2e2e0a00",
  1429 => x"42494f53",
  1430 => x"5f4d3250",
  1431 => x"524f4d00",
  1432 => x"4f70656e",
  1433 => x"65642042",
  1434 => x"494f532c",
  1435 => x"206c6f61",
  1436 => x"64696e67",
  1437 => x"2e2e2e0a",
  1438 => x"00000000",
  1439 => x"52656164",
  1440 => x"20626c6f",
  1441 => x"636b2066",
  1442 => x"61696c65",
  1443 => x"640a0000",
  1444 => x"4c6f6164",
  1445 => x"696e6720",
  1446 => x"42494f53",
  1447 => x"20666169",
  1448 => x"6c65640a",
  1449 => x"00000000",
  1450 => x"52656164",
  1451 => x"206f6620",
  1452 => x"4d425220",
  1453 => x"6661696c",
  1454 => x"65640a00",
  1455 => x"46415431",
  1456 => x"36202020",
  1457 => x"00000000",
  1458 => x"46415433",
  1459 => x"32202020",
  1460 => x"00000000",
  1461 => x"25642070",
  1462 => x"61727469",
  1463 => x"74696f6e",
  1464 => x"7320666f",
  1465 => x"756e640a",
  1466 => x"00000000",
  1467 => x"4e6f2070",
  1468 => x"61727469",
  1469 => x"74696f6e",
  1470 => x"20736967",
  1471 => x"6e617475",
  1472 => x"72652066",
  1473 => x"6f756e64",
  1474 => x"0a000000",
  1475 => x"556e7375",
  1476 => x"70706f72",
  1477 => x"74656420",
  1478 => x"70617274",
  1479 => x"6974696f",
  1480 => x"6e207479",
  1481 => x"7065210a",
  1482 => x"00000000",
  1483 => x"53444843",
  1484 => x"20496e69",
  1485 => x"7469616c",
  1486 => x"697a6174",
  1487 => x"696f6e20",
  1488 => x"6572726f",
  1489 => x"72210a00",
  1490 => x"434d4435",
  1491 => x"38202564",
  1492 => x"0a202000",
  1493 => x"496e6974",
  1494 => x"69616c69",
  1495 => x"73696e67",
  1496 => x"20534420",
  1497 => x"63617264",
  1498 => x"2e2e2e0a",
  1499 => x"00000000",
  1500 => x"53442063",
  1501 => x"61726420",
  1502 => x"72657365",
  1503 => x"74206661",
  1504 => x"696c6564",
  1505 => x"210a0000",
  1506 => x"52656164",
  1507 => x"20636f6d",
  1508 => x"6d616e64",
  1509 => x"20666169",
  1510 => x"6c656420",
  1511 => x"61742025",
  1512 => x"64202825",
  1513 => x"64290a00",
  1514 => x"16200000",
  1515 => x"14200000",
  1516 => x"15200000",
  1517 => x"00000002",
  1518 => x"00000004",
  1519 => x"0000143c",
  1520 => x"000017e8",
  1521 => x"00000002",
  1522 => x"0000144c",
  1523 => x"0000053e",
  1524 => x"00000002",
  1525 => x"00001454",
  1526 => x"0000120b",
  1527 => x"00000000",
  1528 => x"00000000",
  1529 => x"00000000",
  1530 => x"00000003",
  1531 => x"00001878",
  1532 => x"00000003",
  1533 => x"00000001",
  1534 => x"0000145c",
  1535 => x"00000002",
  1536 => x"00000003",
  1537 => x"0000186c",
  1538 => x"00000003",
  1539 => x"00000003",
  1540 => x"0000185c",
  1541 => x"00000004",
  1542 => x"00000001",
  1543 => x"00001464",
  1544 => x"00000006",
  1545 => x"00000001",
  1546 => x"00001480",
  1547 => x"00000007",
  1548 => x"00000003",
  1549 => x"00001854",
  1550 => x"00000002",
  1551 => x"00000004",
  1552 => x"00001494",
  1553 => x"000017b8",
  1554 => x"00000000",
  1555 => x"00000000",
  1556 => x"00000000",
  1557 => x"0000149c",
  1558 => x"000014a8",
  1559 => x"000014b4",
  1560 => x"000014c0",
  1561 => x"000014d8",
  1562 => x"000014f0",
  1563 => x"0000150c",
  1564 => x"00001518",
  1565 => x"00001530",
  1566 => x"00001540",
  1567 => x"00001554",
  1568 => x"00001568",
  1569 => x"00000000",
  1570 => x"00000000",
  1571 => x"00000000",
  1572 => x"00000000",
  1573 => x"00000000",
  1574 => x"00000000",
  1575 => x"00000000",
  1576 => x"00000000",
  1577 => x"00000000",
  1578 => x"00000000",
  1579 => x"00000000",
  1580 => x"00000000",
  1581 => x"00000000",
  1582 => x"00000000",
  1583 => x"00000000",
  1584 => x"00000000",
  1585 => x"00000000",
  1586 => x"00000000",
  1587 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

