-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b0bb7",
     9 => x"ac080b0b",
    10 => x"0bb7b008",
    11 => x"0b0b0bb7",
    12 => x"b4080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"b7b40c0b",
    16 => x"0b0bb7b0",
    17 => x"0c0b0b0b",
    18 => x"b7ac0c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0bae88",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"b7ac70bc",
    57 => x"e4278b38",
    58 => x"80717084",
    59 => x"05530c81",
    60 => x"e2048c51",
    61 => x"8cf40402",
    62 => x"fc050df8",
    63 => x"80518f0b",
    64 => x"b7bc0c9f",
    65 => x"0bb7c00c",
    66 => x"a0717081",
    67 => x"055334b7",
    68 => x"c008ff05",
    69 => x"b7c00cb7",
    70 => x"c0088025",
    71 => x"eb38b7bc",
    72 => x"08ff05b7",
    73 => x"bc0cb7bc",
    74 => x"088025d7",
    75 => x"38028405",
    76 => x"0d0402f0",
    77 => x"050df880",
    78 => x"53f8a054",
    79 => x"83bf5273",
    80 => x"70810555",
    81 => x"33517073",
    82 => x"70810555",
    83 => x"34ff1252",
    84 => x"718025eb",
    85 => x"38fbc053",
    86 => x"9f52a073",
    87 => x"70810555",
    88 => x"34ff1252",
    89 => x"718025f2",
    90 => x"38029005",
    91 => x"0d0402f4",
    92 => x"050d7453",
    93 => x"8e0bb7bc",
    94 => x"08258f38",
    95 => x"82b22db7",
    96 => x"bc08ff05",
    97 => x"b7bc0c82",
    98 => x"f404b7bc",
    99 => x"08b7c008",
   100 => x"5351728a",
   101 => x"2e098106",
   102 => x"b7387151",
   103 => x"719f24a0",
   104 => x"38b7bc08",
   105 => x"a02911f8",
   106 => x"80115151",
   107 => x"a07134b7",
   108 => x"c0088105",
   109 => x"b7c00cb7",
   110 => x"c008519f",
   111 => x"7125e238",
   112 => x"800bb7c0",
   113 => x"0cb7bc08",
   114 => x"8105b7bc",
   115 => x"0c83e404",
   116 => x"70a02912",
   117 => x"f8801151",
   118 => x"51727134",
   119 => x"b7c00881",
   120 => x"05b7c00c",
   121 => x"b7c008a0",
   122 => x"2e098106",
   123 => x"8e38800b",
   124 => x"b7c00cb7",
   125 => x"bc088105",
   126 => x"b7bc0c02",
   127 => x"8c050d04",
   128 => x"02e8050d",
   129 => x"77795656",
   130 => x"880bfc16",
   131 => x"77712c8f",
   132 => x"06545254",
   133 => x"80537272",
   134 => x"25953871",
   135 => x"53fbe014",
   136 => x"51877134",
   137 => x"8114ff14",
   138 => x"545472f1",
   139 => x"387153f9",
   140 => x"1576712c",
   141 => x"87065351",
   142 => x"71802e8b",
   143 => x"38fbe014",
   144 => x"51717134",
   145 => x"81145472",
   146 => x"8e249538",
   147 => x"8f733153",
   148 => x"fbe01451",
   149 => x"a0713481",
   150 => x"14ff1454",
   151 => x"5472f138",
   152 => x"0298050d",
   153 => x"0402ec05",
   154 => x"0d800bb7",
   155 => x"c40cf68c",
   156 => x"08f69008",
   157 => x"71882c56",
   158 => x"5481ff06",
   159 => x"52737225",
   160 => x"88387154",
   161 => x"820bb7c4",
   162 => x"0c72882c",
   163 => x"7381ff06",
   164 => x"54557473",
   165 => x"258b3872",
   166 => x"b7c40884",
   167 => x"07b7c40c",
   168 => x"5573842b",
   169 => x"86a07125",
   170 => x"83713170",
   171 => x"0b0b0bb4",
   172 => x"880c8171",
   173 => x"2bff05f6",
   174 => x"880cfecc",
   175 => x"13ff122c",
   176 => x"788829ff",
   177 => x"94057081",
   178 => x"2cb7c408",
   179 => x"52585255",
   180 => x"51525476",
   181 => x"802e8538",
   182 => x"70810751",
   183 => x"70f6940c",
   184 => x"71098105",
   185 => x"f6800c72",
   186 => x"098105f6",
   187 => x"840c0294",
   188 => x"050d0402",
   189 => x"f4050d74",
   190 => x"53727081",
   191 => x"055480f5",
   192 => x"2d527180",
   193 => x"2e893871",
   194 => x"5182ee2d",
   195 => x"85f90402",
   196 => x"8c050d04",
   197 => x"02f8050d",
   198 => x"a5c12d80",
   199 => x"da51a6f8",
   200 => x"2db7ac08",
   201 => x"812a7081",
   202 => x"06515271",
   203 => x"802ee938",
   204 => x"0288050d",
   205 => x"0402f405",
   206 => x"0dbcd408",
   207 => x"99c406b6",
   208 => x"840b80f5",
   209 => x"2d525270",
   210 => x"802e8638",
   211 => x"71848007",
   212 => x"52b5bc0b",
   213 => x"80f52d72",
   214 => x"07b5e00b",
   215 => x"80f52d70",
   216 => x"812a7081",
   217 => x"06515354",
   218 => x"5270802e",
   219 => x"86387182",
   220 => x"80075272",
   221 => x"81065170",
   222 => x"802e8538",
   223 => x"71880752",
   224 => x"b5ec0b80",
   225 => x"f52d7084",
   226 => x"2b730781",
   227 => x"8432b7ac",
   228 => x"0c51028c",
   229 => x"050d0402",
   230 => x"f4050d74",
   231 => x"70818432",
   232 => x"bcd40c70",
   233 => x"83065253",
   234 => x"70b5b40b",
   235 => x"880581b7",
   236 => x"2d72892a",
   237 => x"70810651",
   238 => x"5170b684",
   239 => x"0b81b72d",
   240 => x"72832a81",
   241 => x"0673882a",
   242 => x"70810651",
   243 => x"52527080",
   244 => x"2e853871",
   245 => x"82075271",
   246 => x"b5e00b81",
   247 => x"b72d7284",
   248 => x"2c708306",
   249 => x"515170b5",
   250 => x"ec0b81b7",
   251 => x"2d70b7ac",
   252 => x"0c028c05",
   253 => x"0d0402f4",
   254 => x"050db4ec",
   255 => x"0b881180",
   256 => x"f52d8c12",
   257 => x"881180f5",
   258 => x"2d70842b",
   259 => x"73078c13",
   260 => x"881180f5",
   261 => x"2d70882b",
   262 => x"73079413",
   263 => x"80f52d70",
   264 => x"8c2b7207",
   265 => x"b7ac0c53",
   266 => x"53535353",
   267 => x"56525351",
   268 => x"028c050d",
   269 => x"0402f405",
   270 => x"0d74b4ec",
   271 => x"71870655",
   272 => x"53517288",
   273 => x"1381b72d",
   274 => x"8c127184",
   275 => x"2c708706",
   276 => x"55525272",
   277 => x"881381b7",
   278 => x"2d8c1271",
   279 => x"842c7087",
   280 => x"06555252",
   281 => x"72881381",
   282 => x"b72d7084",
   283 => x"2c708706",
   284 => x"51517094",
   285 => x"1381b72d",
   286 => x"028c050d",
   287 => x"0402d405",
   288 => x"0db18851",
   289 => x"85f32d9d",
   290 => x"a52db7ac",
   291 => x"08802e83",
   292 => x"893886b5",
   293 => x"2db7ac08",
   294 => x"538fee2d",
   295 => x"b7ac0854",
   296 => x"b7ac0880",
   297 => x"2e82f538",
   298 => x"a1a82db7",
   299 => x"ac08802e",
   300 => x"8738b1a0",
   301 => x"5189c504",
   302 => x"99912db7",
   303 => x"ac08802e",
   304 => x"a238b1b4",
   305 => x"5185f32d",
   306 => x"b1cc5185",
   307 => x"f32d8694",
   308 => x"2d728407",
   309 => x"53810bfe",
   310 => x"c40c72fe",
   311 => x"c00c7251",
   312 => x"87972d84",
   313 => x"0bfec40c",
   314 => x"7c802eab",
   315 => x"38b1e852",
   316 => x"b7cc5196",
   317 => x"802db7ac",
   318 => x"08802e80",
   319 => x"c33872b7",
   320 => x"d80c87f6",
   321 => x"2db7ac08",
   322 => x"b7dc0cb7",
   323 => x"d852b7cc",
   324 => x"5198eb2d",
   325 => x"8ac004b1",
   326 => x"e852b7cc",
   327 => x"5196802d",
   328 => x"b7ac0880",
   329 => x"2e9a38b7",
   330 => x"d852b7cc",
   331 => x"5198c52d",
   332 => x"b7d808b7",
   333 => x"dc085253",
   334 => x"88b52d72",
   335 => x"5187972d",
   336 => x"b1f45185",
   337 => x"f32db28c",
   338 => x"52b7cc51",
   339 => x"96802db7",
   340 => x"ac089838",
   341 => x"b2985185",
   342 => x"f32db2b0",
   343 => x"52b7cc51",
   344 => x"96802db7",
   345 => x"ac08802e",
   346 => x"81b038b2",
   347 => x"bc5185f3",
   348 => x"2db7d008",
   349 => x"57807759",
   350 => x"5a767a2e",
   351 => x"8b38811a",
   352 => x"78812a59",
   353 => x"5a77f738",
   354 => x"f71a5a80",
   355 => x"77258180",
   356 => x"38795277",
   357 => x"5184802d",
   358 => x"b7d852b7",
   359 => x"cc5198c5",
   360 => x"2db7ac08",
   361 => x"53b7ac08",
   362 => x"802e80c9",
   363 => x"38b7d85b",
   364 => x"80598be2",
   365 => x"047a7084",
   366 => x"055c0870",
   367 => x"81ff0671",
   368 => x"882c7081",
   369 => x"ff067390",
   370 => x"2c7081ff",
   371 => x"0675982a",
   372 => x"fec80cfe",
   373 => x"c80c58fe",
   374 => x"c80c57fe",
   375 => x"c80c841a",
   376 => x"5a537653",
   377 => x"84807725",
   378 => x"84388480",
   379 => x"53727924",
   380 => x"c4388c80",
   381 => x"04b2cc51",
   382 => x"85f32d72",
   383 => x"548c9c04",
   384 => x"b7cc5198",
   385 => x"982dfc80",
   386 => x"17811959",
   387 => x"578b8b04",
   388 => x"820bfec4",
   389 => x"0c81548c",
   390 => x"9c048054",
   391 => x"73b7ac0c",
   392 => x"02ac050d",
   393 => x"0402f805",
   394 => x"0da7c82d",
   395 => x"81f72d81",
   396 => x"5184e52d",
   397 => x"fec45281",
   398 => x"720ca588",
   399 => x"2da5882d",
   400 => x"84720c73",
   401 => x"5188fd2d",
   402 => x"b48c51a9",
   403 => x"a62d8051",
   404 => x"84e52d02",
   405 => x"88050d04",
   406 => x"02fc050d",
   407 => x"81518ca5",
   408 => x"2d028405",
   409 => x"0d0402fc",
   410 => x"050d8051",
   411 => x"8ca52d02",
   412 => x"84050d04",
   413 => x"02ec050d",
   414 => x"8cb85187",
   415 => x"972d810b",
   416 => x"fec40c8c",
   417 => x"b80bfec0",
   418 => x"0c840bfe",
   419 => x"c40c830b",
   420 => x"fecc0ca5",
   421 => x"a32da7bc",
   422 => x"2da5882d",
   423 => x"a5882d81",
   424 => x"f72d8151",
   425 => x"84e52da5",
   426 => x"882da588",
   427 => x"2d815184",
   428 => x"e52d8051",
   429 => x"88fd2db7",
   430 => x"ac08802e",
   431 => x"81dd3880",
   432 => x"5184e52d",
   433 => x"b48c51a9",
   434 => x"a62dbcbc",
   435 => x"08097083",
   436 => x"06fecc0c",
   437 => x"52bcb408",
   438 => x"8938bcb8",
   439 => x"08802e80",
   440 => x"e238fed0",
   441 => x"08708106",
   442 => x"51527180",
   443 => x"2e80d438",
   444 => x"a7c22dbc",
   445 => x"b40870bc",
   446 => x"b8087057",
   447 => x"55565280",
   448 => x"ff722584",
   449 => x"3880ff52",
   450 => x"80ff7325",
   451 => x"843880ff",
   452 => x"5371ff80",
   453 => x"258438ff",
   454 => x"805272ff",
   455 => x"80258438",
   456 => x"ff805374",
   457 => x"7231bcb4",
   458 => x"0c737331",
   459 => x"bcb80ca7",
   460 => x"bc2d7188",
   461 => x"2b83fe80",
   462 => x"067381ff",
   463 => x"067107fe",
   464 => x"d00c52a5",
   465 => x"c12da9b6",
   466 => x"2db7ac08",
   467 => x"5386b52d",
   468 => x"b7ac08fe",
   469 => x"c00c87f6",
   470 => x"2db7ac08",
   471 => x"fed40c86",
   472 => x"b52db7ac",
   473 => x"08b7c808",
   474 => x"2e9c38b7",
   475 => x"ac08b7c8",
   476 => x"0c845272",
   477 => x"5184e52d",
   478 => x"a5882da5",
   479 => x"882dff12",
   480 => x"52718025",
   481 => x"ee387280",
   482 => x"2e89388a",
   483 => x"0bfec40c",
   484 => x"8dca0482",
   485 => x"0bfec40c",
   486 => x"8dca04b2",
   487 => x"dc5185f3",
   488 => x"2d820bfe",
   489 => x"c40c800b",
   490 => x"b7ac0c02",
   491 => x"94050d04",
   492 => x"02e8050d",
   493 => x"77797b58",
   494 => x"55558053",
   495 => x"727625a3",
   496 => x"38747081",
   497 => x"055680f5",
   498 => x"2d747081",
   499 => x"055680f5",
   500 => x"2d525271",
   501 => x"712e8638",
   502 => x"81518fe5",
   503 => x"04811353",
   504 => x"8fbc0480",
   505 => x"5170b7ac",
   506 => x"0c029805",
   507 => x"0d0402d8",
   508 => x"050d800b",
   509 => x"bbe00cb7",
   510 => x"d8528051",
   511 => x"a08d2db7",
   512 => x"ac0854b7",
   513 => x"ac088c38",
   514 => x"b2f45185",
   515 => x"f32d7355",
   516 => x"95890480",
   517 => x"56810bbc",
   518 => x"840c8853",
   519 => x"b38052b8",
   520 => x"8e518fb0",
   521 => x"2db7ac08",
   522 => x"762e0981",
   523 => x"068738b7",
   524 => x"ac08bc84",
   525 => x"0c8853b3",
   526 => x"8c52b8aa",
   527 => x"518fb02d",
   528 => x"b7ac0887",
   529 => x"38b7ac08",
   530 => x"bc840cbc",
   531 => x"8408802e",
   532 => x"80f638bb",
   533 => x"9e0b80f5",
   534 => x"2dbb9f0b",
   535 => x"80f52d71",
   536 => x"982b7190",
   537 => x"2b07bba0",
   538 => x"0b80f52d",
   539 => x"70882b72",
   540 => x"07bba10b",
   541 => x"80f52d71",
   542 => x"07bbd60b",
   543 => x"80f52dbb",
   544 => x"d70b80f5",
   545 => x"2d71882b",
   546 => x"07535f54",
   547 => x"525a5657",
   548 => x"557381ab",
   549 => x"aa2e0981",
   550 => x"068d3875",
   551 => x"51a1af2d",
   552 => x"b7ac0856",
   553 => x"91b40473",
   554 => x"82d4d52e",
   555 => x"8738b398",
   556 => x"5191f504",
   557 => x"b7d85275",
   558 => x"51a08d2d",
   559 => x"b7ac0855",
   560 => x"b7ac0880",
   561 => x"2e83c238",
   562 => x"8853b38c",
   563 => x"52b8aa51",
   564 => x"8fb02db7",
   565 => x"ac088938",
   566 => x"810bbbe0",
   567 => x"0c91fb04",
   568 => x"8853b380",
   569 => x"52b88e51",
   570 => x"8fb02db7",
   571 => x"ac08802e",
   572 => x"8a38b3ac",
   573 => x"5185f32d",
   574 => x"92d504bb",
   575 => x"d60b80f5",
   576 => x"2d547380",
   577 => x"d52e0981",
   578 => x"0680ca38",
   579 => x"bbd70b80",
   580 => x"f52d5473",
   581 => x"81aa2e09",
   582 => x"8106ba38",
   583 => x"800bb7d8",
   584 => x"0b80f52d",
   585 => x"56547481",
   586 => x"e92e8338",
   587 => x"81547481",
   588 => x"eb2e8c38",
   589 => x"80557375",
   590 => x"2e098106",
   591 => x"82cb38b7",
   592 => x"e30b80f5",
   593 => x"2d55748d",
   594 => x"38b7e40b",
   595 => x"80f52d54",
   596 => x"73822e86",
   597 => x"38805595",
   598 => x"8904b7e5",
   599 => x"0b80f52d",
   600 => x"70bbd80c",
   601 => x"ff05bbdc",
   602 => x"0cb7e60b",
   603 => x"80f52db7",
   604 => x"e70b80f5",
   605 => x"2d587605",
   606 => x"77828029",
   607 => x"0570bbe4",
   608 => x"0cb7e80b",
   609 => x"80f52d70",
   610 => x"bbf80cbb",
   611 => x"e0085957",
   612 => x"5876802e",
   613 => x"81a33888",
   614 => x"53b38c52",
   615 => x"b8aa518f",
   616 => x"b02db7ac",
   617 => x"0881e238",
   618 => x"bbd80870",
   619 => x"842bbbfc",
   620 => x"0c70bbf4",
   621 => x"0cb7fd0b",
   622 => x"80f52db7",
   623 => x"fc0b80f5",
   624 => x"2d718280",
   625 => x"2905b7fe",
   626 => x"0b80f52d",
   627 => x"70848080",
   628 => x"2912b7ff",
   629 => x"0b80f52d",
   630 => x"7081800a",
   631 => x"291270bc",
   632 => x"800cbbf8",
   633 => x"087129bb",
   634 => x"e4080570",
   635 => x"bbe80cb8",
   636 => x"850b80f5",
   637 => x"2db8840b",
   638 => x"80f52d71",
   639 => x"82802905",
   640 => x"b8860b80",
   641 => x"f52d7084",
   642 => x"80802912",
   643 => x"b8870b80",
   644 => x"f52d7098",
   645 => x"2b81f00a",
   646 => x"06720570",
   647 => x"bbec0cfe",
   648 => x"117e2977",
   649 => x"05bbf00c",
   650 => x"52595243",
   651 => x"545e5152",
   652 => x"59525d57",
   653 => x"59579587",
   654 => x"04b7ea0b",
   655 => x"80f52db7",
   656 => x"e90b80f5",
   657 => x"2d718280",
   658 => x"290570bb",
   659 => x"fc0c70a0",
   660 => x"2983ff05",
   661 => x"70892a70",
   662 => x"bbf40cb7",
   663 => x"ef0b80f5",
   664 => x"2db7ee0b",
   665 => x"80f52d71",
   666 => x"82802905",
   667 => x"70bc800c",
   668 => x"7b71291e",
   669 => x"70bbf00c",
   670 => x"7dbbec0c",
   671 => x"7305bbe8",
   672 => x"0c555e51",
   673 => x"51555581",
   674 => x"5574b7ac",
   675 => x"0c02a805",
   676 => x"0d0402ec",
   677 => x"050d7670",
   678 => x"872c7180",
   679 => x"ff065556",
   680 => x"54bbe008",
   681 => x"8a387388",
   682 => x"2c7481ff",
   683 => x"065455b7",
   684 => x"d852bbe4",
   685 => x"081551a0",
   686 => x"8d2db7ac",
   687 => x"0854b7ac",
   688 => x"08802eb3",
   689 => x"38bbe008",
   690 => x"802e9838",
   691 => x"728429b7",
   692 => x"d8057008",
   693 => x"5253a1af",
   694 => x"2db7ac08",
   695 => x"f00a0653",
   696 => x"95f50472",
   697 => x"10b7d805",
   698 => x"7080e02d",
   699 => x"5253a1df",
   700 => x"2db7ac08",
   701 => x"53725473",
   702 => x"b7ac0c02",
   703 => x"94050d04",
   704 => x"02c8050d",
   705 => x"7f615f5b",
   706 => x"800bbbec",
   707 => x"08bbf008",
   708 => x"595d56bb",
   709 => x"e008762e",
   710 => x"8a38bbd8",
   711 => x"08842b58",
   712 => x"96a904bb",
   713 => x"f408842b",
   714 => x"58805978",
   715 => x"782781a9",
   716 => x"38788f06",
   717 => x"a0175754",
   718 => x"738f38b7",
   719 => x"d8527651",
   720 => x"811757a0",
   721 => x"8d2db7d8",
   722 => x"56807680",
   723 => x"f52d5654",
   724 => x"74742e83",
   725 => x"38815474",
   726 => x"81e52e80",
   727 => x"f6388170",
   728 => x"7506555d",
   729 => x"73802e80",
   730 => x"ea388b16",
   731 => x"80f52d98",
   732 => x"065a7980",
   733 => x"de388b53",
   734 => x"7d527551",
   735 => x"8fb02db7",
   736 => x"ac0880cf",
   737 => x"389c1608",
   738 => x"51a1af2d",
   739 => x"b7ac0884",
   740 => x"1c0c9a16",
   741 => x"80e02d51",
   742 => x"a1df2db7",
   743 => x"ac08b7ac",
   744 => x"08881d0c",
   745 => x"b7ac0855",
   746 => x"55bbe008",
   747 => x"802e9838",
   748 => x"941680e0",
   749 => x"2d51a1df",
   750 => x"2db7ac08",
   751 => x"902b83ff",
   752 => x"f00a0670",
   753 => x"16515473",
   754 => x"881c0c79",
   755 => x"7b0c7c54",
   756 => x"988f0481",
   757 => x"195996ab",
   758 => x"04bbe008",
   759 => x"802eae38",
   760 => x"7b519592",
   761 => x"2db7ac08",
   762 => x"b7ac0880",
   763 => x"fffffff8",
   764 => x"06555c73",
   765 => x"80ffffff",
   766 => x"f82e9238",
   767 => x"b7ac08fe",
   768 => x"05bbd808",
   769 => x"29bbe808",
   770 => x"055796a9",
   771 => x"04805473",
   772 => x"b7ac0c02",
   773 => x"b8050d04",
   774 => x"02f4050d",
   775 => x"74700881",
   776 => x"05710c70",
   777 => x"08bbdc08",
   778 => x"06535371",
   779 => x"8e388813",
   780 => x"08519592",
   781 => x"2db7ac08",
   782 => x"88140c81",
   783 => x"0bb7ac0c",
   784 => x"028c050d",
   785 => x"0402f005",
   786 => x"0d758811",
   787 => x"08fe05bb",
   788 => x"d80829bb",
   789 => x"e8081172",
   790 => x"08bbdc08",
   791 => x"06057955",
   792 => x"535454a0",
   793 => x"8d2d0290",
   794 => x"050d0402",
   795 => x"f0050d75",
   796 => x"881108fe",
   797 => x"05bbd808",
   798 => x"29bbe808",
   799 => x"117208bb",
   800 => x"dc080605",
   801 => x"79555354",
   802 => x"549ecd2d",
   803 => x"0290050d",
   804 => x"04bbe008",
   805 => x"b7ac0c04",
   806 => x"02f4050d",
   807 => x"d45281ff",
   808 => x"720c7108",
   809 => x"5381ff72",
   810 => x"0c72882b",
   811 => x"83fe8006",
   812 => x"72087081",
   813 => x"ff065152",
   814 => x"5381ff72",
   815 => x"0c727107",
   816 => x"882b7208",
   817 => x"7081ff06",
   818 => x"51525381",
   819 => x"ff720c72",
   820 => x"7107882b",
   821 => x"72087081",
   822 => x"ff067207",
   823 => x"b7ac0c52",
   824 => x"53028c05",
   825 => x"0d0402f4",
   826 => x"050d7476",
   827 => x"7181ff06",
   828 => x"d40c5353",
   829 => x"bc880885",
   830 => x"3871892b",
   831 => x"5271982a",
   832 => x"d40c7190",
   833 => x"2a7081ff",
   834 => x"06d40c51",
   835 => x"71882a70",
   836 => x"81ff06d4",
   837 => x"0c517181",
   838 => x"ff06d40c",
   839 => x"72902a70",
   840 => x"81ff06d4",
   841 => x"0c51d408",
   842 => x"7081ff06",
   843 => x"515182b8",
   844 => x"bf527081",
   845 => x"ff2e0981",
   846 => x"06943881",
   847 => x"ff0bd40c",
   848 => x"d4087081",
   849 => x"ff06ff14",
   850 => x"54515171",
   851 => x"e53870b7",
   852 => x"ac0c028c",
   853 => x"050d0402",
   854 => x"fc050d81",
   855 => x"c75181ff",
   856 => x"0bd40cff",
   857 => x"11517080",
   858 => x"25f43802",
   859 => x"84050d04",
   860 => x"02f0050d",
   861 => x"9ad72d8f",
   862 => x"cf538052",
   863 => x"87fc80f7",
   864 => x"5199e62d",
   865 => x"b7ac0854",
   866 => x"b7ac0881",
   867 => x"2e098106",
   868 => x"a33881ff",
   869 => x"0bd40c82",
   870 => x"0a52849c",
   871 => x"80e95199",
   872 => x"e62db7ac",
   873 => x"088b3881",
   874 => x"ff0bd40c",
   875 => x"73539bba",
   876 => x"049ad72d",
   877 => x"ff135372",
   878 => x"c13872b7",
   879 => x"ac0c0290",
   880 => x"050d0402",
   881 => x"f4050d81",
   882 => x"ff0bd40c",
   883 => x"93538052",
   884 => x"87fc80c1",
   885 => x"5199e62d",
   886 => x"b7ac088b",
   887 => x"3881ff0b",
   888 => x"d40c8153",
   889 => x"9bf0049a",
   890 => x"d72dff13",
   891 => x"5372df38",
   892 => x"72b7ac0c",
   893 => x"028c050d",
   894 => x"0402f005",
   895 => x"0d9ad72d",
   896 => x"83aa5284",
   897 => x"9c80c851",
   898 => x"99e62db7",
   899 => x"ac08812e",
   900 => x"09810692",
   901 => x"3899982d",
   902 => x"b7ac0883",
   903 => x"ffff0653",
   904 => x"7283aa2e",
   905 => x"97389bc3",
   906 => x"2d9cb704",
   907 => x"81549d9c",
   908 => x"04b3b851",
   909 => x"85f32d80",
   910 => x"549d9c04",
   911 => x"81ff0bd4",
   912 => x"0cb1539a",
   913 => x"f02db7ac",
   914 => x"08802e80",
   915 => x"c0388052",
   916 => x"87fc80fa",
   917 => x"5199e62d",
   918 => x"b7ac08b1",
   919 => x"3881ff0b",
   920 => x"d40cd408",
   921 => x"5381ff0b",
   922 => x"d40c81ff",
   923 => x"0bd40c81",
   924 => x"ff0bd40c",
   925 => x"81ff0bd4",
   926 => x"0c72862a",
   927 => x"708106b7",
   928 => x"ac085651",
   929 => x"5372802e",
   930 => x"93389cac",
   931 => x"0472822e",
   932 => x"ff9f38ff",
   933 => x"135372ff",
   934 => x"aa387254",
   935 => x"73b7ac0c",
   936 => x"0290050d",
   937 => x"0402f005",
   938 => x"0d810bbc",
   939 => x"880c8454",
   940 => x"d008708f",
   941 => x"2a708106",
   942 => x"51515372",
   943 => x"f33872d0",
   944 => x"0c9ad72d",
   945 => x"b3c85185",
   946 => x"f32dd008",
   947 => x"708f2a70",
   948 => x"81065151",
   949 => x"5372f338",
   950 => x"810bd00c",
   951 => x"b1538052",
   952 => x"84d480c0",
   953 => x"5199e62d",
   954 => x"b7ac0881",
   955 => x"2ea13872",
   956 => x"822e0981",
   957 => x"068c38b3",
   958 => x"d45185f3",
   959 => x"2d80539e",
   960 => x"c404ff13",
   961 => x"5372d738",
   962 => x"ff145473",
   963 => x"ffa2389b",
   964 => x"f92db7ac",
   965 => x"08bc880c",
   966 => x"b7ac088b",
   967 => x"38815287",
   968 => x"fc80d051",
   969 => x"99e62d81",
   970 => x"ff0bd40c",
   971 => x"d008708f",
   972 => x"2a708106",
   973 => x"51515372",
   974 => x"f33872d0",
   975 => x"0c81ff0b",
   976 => x"d40c8153",
   977 => x"72b7ac0c",
   978 => x"0290050d",
   979 => x"0402e805",
   980 => x"0d785681",
   981 => x"ff0bd40c",
   982 => x"d008708f",
   983 => x"2a708106",
   984 => x"51515372",
   985 => x"f3388281",
   986 => x"0bd00c81",
   987 => x"ff0bd40c",
   988 => x"775287fc",
   989 => x"80d85199",
   990 => x"e62db7ac",
   991 => x"08802e8c",
   992 => x"38b3ec51",
   993 => x"85f32d81",
   994 => x"53a08404",
   995 => x"81ff0bd4",
   996 => x"0c81fe0b",
   997 => x"d40c80ff",
   998 => x"55757084",
   999 => x"05570870",
  1000 => x"982ad40c",
  1001 => x"70902c70",
  1002 => x"81ff06d4",
  1003 => x"0c547088",
  1004 => x"2c7081ff",
  1005 => x"06d40c54",
  1006 => x"7081ff06",
  1007 => x"d40c54ff",
  1008 => x"15557480",
  1009 => x"25d33881",
  1010 => x"ff0bd40c",
  1011 => x"81ff0bd4",
  1012 => x"0c81ff0b",
  1013 => x"d40c868d",
  1014 => x"a05481ff",
  1015 => x"0bd40cd4",
  1016 => x"0881ff06",
  1017 => x"55748738",
  1018 => x"ff145473",
  1019 => x"ed3881ff",
  1020 => x"0bd40cd0",
  1021 => x"08708f2a",
  1022 => x"70810651",
  1023 => x"515372f3",
  1024 => x"3872d00c",
  1025 => x"72b7ac0c",
  1026 => x"0298050d",
  1027 => x"0402e805",
  1028 => x"0d785580",
  1029 => x"5681ff0b",
  1030 => x"d40cd008",
  1031 => x"708f2a70",
  1032 => x"81065151",
  1033 => x"5372f338",
  1034 => x"82810bd0",
  1035 => x"0c81ff0b",
  1036 => x"d40c7752",
  1037 => x"87fc80d1",
  1038 => x"5199e62d",
  1039 => x"80dbc6df",
  1040 => x"54b7ac08",
  1041 => x"802e8a38",
  1042 => x"b2cc5185",
  1043 => x"f32da19f",
  1044 => x"0481ff0b",
  1045 => x"d40cd408",
  1046 => x"7081ff06",
  1047 => x"51537281",
  1048 => x"fe2e0981",
  1049 => x"069d3880",
  1050 => x"ff539998",
  1051 => x"2db7ac08",
  1052 => x"75708405",
  1053 => x"570cff13",
  1054 => x"53728025",
  1055 => x"ed388156",
  1056 => x"a18904ff",
  1057 => x"145473c9",
  1058 => x"3881ff0b",
  1059 => x"d40cd008",
  1060 => x"708f2a70",
  1061 => x"81065151",
  1062 => x"5372f338",
  1063 => x"72d00c75",
  1064 => x"b7ac0c02",
  1065 => x"98050d04",
  1066 => x"bc8808b7",
  1067 => x"ac0c0402",
  1068 => x"f4050d74",
  1069 => x"70882a83",
  1070 => x"fe800670",
  1071 => x"72982a07",
  1072 => x"72882b87",
  1073 => x"fc808006",
  1074 => x"73982b81",
  1075 => x"f00a0671",
  1076 => x"730707b7",
  1077 => x"ac0c5651",
  1078 => x"5351028c",
  1079 => x"050d0402",
  1080 => x"f8050d02",
  1081 => x"8e0580f5",
  1082 => x"2d74882b",
  1083 => x"077083ff",
  1084 => x"ff06b7ac",
  1085 => x"0c510288",
  1086 => x"050d0402",
  1087 => x"fc050d72",
  1088 => x"5180710c",
  1089 => x"800b8412",
  1090 => x"0c028405",
  1091 => x"0d0402f0",
  1092 => x"050d7570",
  1093 => x"08841208",
  1094 => x"535353ff",
  1095 => x"5471712e",
  1096 => x"a838a7c2",
  1097 => x"2d841308",
  1098 => x"70842914",
  1099 => x"88117008",
  1100 => x"7081ff06",
  1101 => x"84180881",
  1102 => x"11870684",
  1103 => x"1a0c5351",
  1104 => x"55515151",
  1105 => x"a7bc2d71",
  1106 => x"5473b7ac",
  1107 => x"0c029005",
  1108 => x"0d0402f0",
  1109 => x"050da7c2",
  1110 => x"2de008e4",
  1111 => x"08718b2a",
  1112 => x"70810651",
  1113 => x"53555270",
  1114 => x"802e9d38",
  1115 => x"bc8c0870",
  1116 => x"8429bc94",
  1117 => x"057381ff",
  1118 => x"06710c51",
  1119 => x"51bc8c08",
  1120 => x"81118706",
  1121 => x"bc8c0c51",
  1122 => x"738b2a70",
  1123 => x"81065151",
  1124 => x"70802e81",
  1125 => x"8938b6dc",
  1126 => x"088429bc",
  1127 => x"c4057481",
  1128 => x"ff06710c",
  1129 => x"51b6dc08",
  1130 => x"8105b6dc",
  1131 => x"0c850bb6",
  1132 => x"d80cb6dc",
  1133 => x"08b6d408",
  1134 => x"2e098106",
  1135 => x"81863880",
  1136 => x"0bb6dc0c",
  1137 => x"bcc40870",
  1138 => x"8306bcbc",
  1139 => x"0c70852a",
  1140 => x"708106bc",
  1141 => x"b8085651",
  1142 => x"52527080",
  1143 => x"2e8e38bc",
  1144 => x"cc08fe80",
  1145 => x"3213bcb8",
  1146 => x"0ca3f304",
  1147 => x"bccc0813",
  1148 => x"bcb80c71",
  1149 => x"842a7081",
  1150 => x"06bcb408",
  1151 => x"54515170",
  1152 => x"802e9038",
  1153 => x"bcc80881",
  1154 => x"ff321281",
  1155 => x"05bcb40c",
  1156 => x"a4c40471",
  1157 => x"bcc80831",
  1158 => x"bcb40ca4",
  1159 => x"c404b6d8",
  1160 => x"08ff05b6",
  1161 => x"d80cb6d8",
  1162 => x"08ff2e09",
  1163 => x"81069538",
  1164 => x"b6dc0880",
  1165 => x"2e8a3887",
  1166 => x"0bb6d408",
  1167 => x"31b6d40c",
  1168 => x"70b6dc0c",
  1169 => x"738a2a70",
  1170 => x"81065151",
  1171 => x"70802e92",
  1172 => x"38b6d008",
  1173 => x"51ff7125",
  1174 => x"893870e4",
  1175 => x"0cff0bb6",
  1176 => x"d00c800b",
  1177 => x"bcc00ca7",
  1178 => x"b52da7bc",
  1179 => x"2d029005",
  1180 => x"0d0402fc",
  1181 => x"050db6d0",
  1182 => x"08517080",
  1183 => x"24fc3872",
  1184 => x"b6d00c02",
  1185 => x"84050d04",
  1186 => x"02fc050d",
  1187 => x"a7c22d81",
  1188 => x"0bbcc00c",
  1189 => x"a7bc2dbc",
  1190 => x"c0085170",
  1191 => x"fa380284",
  1192 => x"050d0402",
  1193 => x"fc050dbc",
  1194 => x"8c51a1fb",
  1195 => x"2da2d251",
  1196 => x"a7b12da6",
  1197 => x"db2d81f4",
  1198 => x"51a4f22d",
  1199 => x"0284050d",
  1200 => x"0402f405",
  1201 => x"0da6c304",
  1202 => x"b7ac0881",
  1203 => x"f02e0981",
  1204 => x"06893881",
  1205 => x"0bb7a00c",
  1206 => x"a6c304b7",
  1207 => x"ac0881e0",
  1208 => x"2e098106",
  1209 => x"8938810b",
  1210 => x"b7a40ca6",
  1211 => x"c304b7ac",
  1212 => x"0852b7a4",
  1213 => x"08802e88",
  1214 => x"38b7ac08",
  1215 => x"81800552",
  1216 => x"71842c72",
  1217 => x"8f065353",
  1218 => x"b7a00880",
  1219 => x"2e993872",
  1220 => x"8429b6e0",
  1221 => x"05721381",
  1222 => x"712b7009",
  1223 => x"73080673",
  1224 => x"0c515353",
  1225 => x"a6b90472",
  1226 => x"8429b6e0",
  1227 => x"05721383",
  1228 => x"712b7208",
  1229 => x"07720c53",
  1230 => x"53800bb7",
  1231 => x"a40c800b",
  1232 => x"b7a00cbc",
  1233 => x"8c51a28e",
  1234 => x"2db7ac08",
  1235 => x"ff24fef8",
  1236 => x"38800bb7",
  1237 => x"ac0c028c",
  1238 => x"050d0402",
  1239 => x"f8050db6",
  1240 => x"e0528f51",
  1241 => x"80727084",
  1242 => x"05540cff",
  1243 => x"11517080",
  1244 => x"25f23802",
  1245 => x"88050d04",
  1246 => x"02f0050d",
  1247 => x"7551a7c2",
  1248 => x"2d70822c",
  1249 => x"fc06b6e0",
  1250 => x"1172109e",
  1251 => x"06710870",
  1252 => x"722a7083",
  1253 => x"0682742b",
  1254 => x"70097406",
  1255 => x"760c5451",
  1256 => x"56575351",
  1257 => x"53a7bc2d",
  1258 => x"71b7ac0c",
  1259 => x"0290050d",
  1260 => x"0471980c",
  1261 => x"04ffb008",
  1262 => x"b7ac0c04",
  1263 => x"810bffb0",
  1264 => x"0c04800b",
  1265 => x"ffb00c04",
  1266 => x"02fc050d",
  1267 => x"800bb7a8",
  1268 => x"0c805184",
  1269 => x"e52d0284",
  1270 => x"050d0402",
  1271 => x"ec050d76",
  1272 => x"54805287",
  1273 => x"0b881580",
  1274 => x"f52d5653",
  1275 => x"74722483",
  1276 => x"38a05372",
  1277 => x"5182ee2d",
  1278 => x"81128b15",
  1279 => x"80f52d54",
  1280 => x"52727225",
  1281 => x"de380294",
  1282 => x"050d0402",
  1283 => x"f0050dbc",
  1284 => x"d8085481",
  1285 => x"f72d800b",
  1286 => x"bcdc0c73",
  1287 => x"08802e81",
  1288 => x"8038820b",
  1289 => x"b7c00cbc",
  1290 => x"dc088f06",
  1291 => x"b7bc0c73",
  1292 => x"08527183",
  1293 => x"2e963871",
  1294 => x"83268938",
  1295 => x"71812eaf",
  1296 => x"38a98c04",
  1297 => x"71852e9f",
  1298 => x"38a98c04",
  1299 => x"881480f5",
  1300 => x"2d841508",
  1301 => x"b3fc5354",
  1302 => x"5285f32d",
  1303 => x"71842913",
  1304 => x"70085252",
  1305 => x"a9900473",
  1306 => x"51a7db2d",
  1307 => x"a98c04bc",
  1308 => x"d4088815",
  1309 => x"082c7081",
  1310 => x"06515271",
  1311 => x"802e8738",
  1312 => x"b48051a9",
  1313 => x"8904b484",
  1314 => x"5185f32d",
  1315 => x"84140851",
  1316 => x"85f32dbc",
  1317 => x"dc088105",
  1318 => x"bcdc0c8c",
  1319 => x"1454a89b",
  1320 => x"04029005",
  1321 => x"0d0471bc",
  1322 => x"d80ca88b",
  1323 => x"2dbcdc08",
  1324 => x"ff05bce0",
  1325 => x"0c0402ec",
  1326 => x"050dbcd8",
  1327 => x"085580f8",
  1328 => x"51a6f82d",
  1329 => x"b7ac0881",
  1330 => x"2a708106",
  1331 => x"5152719b",
  1332 => x"388751a6",
  1333 => x"f82db7ac",
  1334 => x"08812a70",
  1335 => x"81065152",
  1336 => x"71802eb1",
  1337 => x"38a9eb04",
  1338 => x"a5c12d87",
  1339 => x"51a6f82d",
  1340 => x"b7ac08f4",
  1341 => x"38a9fb04",
  1342 => x"a5c12d80",
  1343 => x"f851a6f8",
  1344 => x"2db7ac08",
  1345 => x"f338b7a8",
  1346 => x"08813270",
  1347 => x"b7a80c70",
  1348 => x"525284e5",
  1349 => x"2db7a808",
  1350 => x"a23880da",
  1351 => x"51a6f82d",
  1352 => x"81f551a6",
  1353 => x"f82d81f2",
  1354 => x"51a6f82d",
  1355 => x"81eb51a6",
  1356 => x"f82d81f4",
  1357 => x"51a6f82d",
  1358 => x"adff0481",
  1359 => x"f551a6f8",
  1360 => x"2db7ac08",
  1361 => x"812a7081",
  1362 => x"06515271",
  1363 => x"802e8f38",
  1364 => x"bce00852",
  1365 => x"71802e86",
  1366 => x"38ff12bc",
  1367 => x"e00c81f2",
  1368 => x"51a6f82d",
  1369 => x"b7ac0881",
  1370 => x"2a708106",
  1371 => x"51527180",
  1372 => x"2e9538bc",
  1373 => x"dc08ff05",
  1374 => x"bce00854",
  1375 => x"52727225",
  1376 => x"86388113",
  1377 => x"bce00cbc",
  1378 => x"e0087053",
  1379 => x"5473802e",
  1380 => x"8a388c15",
  1381 => x"ff155555",
  1382 => x"ab8d0482",
  1383 => x"0bb7c00c",
  1384 => x"718f06b7",
  1385 => x"bc0c81eb",
  1386 => x"51a6f82d",
  1387 => x"b7ac0881",
  1388 => x"2a708106",
  1389 => x"51527180",
  1390 => x"2ead3874",
  1391 => x"08852e09",
  1392 => x"8106a438",
  1393 => x"881580f5",
  1394 => x"2dff0552",
  1395 => x"71881681",
  1396 => x"b72d7198",
  1397 => x"2b527180",
  1398 => x"25883880",
  1399 => x"0b881681",
  1400 => x"b72d7451",
  1401 => x"a7db2d81",
  1402 => x"f451a6f8",
  1403 => x"2db7ac08",
  1404 => x"812a7081",
  1405 => x"06515271",
  1406 => x"802eb338",
  1407 => x"7408852e",
  1408 => x"098106aa",
  1409 => x"38881580",
  1410 => x"f52d8105",
  1411 => x"52718816",
  1412 => x"81b72d71",
  1413 => x"81ff068b",
  1414 => x"1680f52d",
  1415 => x"54527272",
  1416 => x"27873872",
  1417 => x"881681b7",
  1418 => x"2d7451a7",
  1419 => x"db2d80da",
  1420 => x"51a6f82d",
  1421 => x"b7ac0881",
  1422 => x"2a708106",
  1423 => x"51527180",
  1424 => x"2e80fb38",
  1425 => x"bcd808bc",
  1426 => x"e0085553",
  1427 => x"73802e8a",
  1428 => x"388c13ff",
  1429 => x"155553ac",
  1430 => x"cc047208",
  1431 => x"5271822e",
  1432 => x"a6387182",
  1433 => x"26893871",
  1434 => x"812ea538",
  1435 => x"adbe0471",
  1436 => x"832ead38",
  1437 => x"71842e09",
  1438 => x"810680c2",
  1439 => x"38881308",
  1440 => x"51a9a62d",
  1441 => x"adbe0488",
  1442 => x"13085271",
  1443 => x"2dadbe04",
  1444 => x"810b8814",
  1445 => x"082bbcd4",
  1446 => x"0832bcd4",
  1447 => x"0cadbb04",
  1448 => x"881380f5",
  1449 => x"2d81058b",
  1450 => x"1480f52d",
  1451 => x"53547174",
  1452 => x"24833880",
  1453 => x"54738814",
  1454 => x"81b72da8",
  1455 => x"8b2d8054",
  1456 => x"800bb7c0",
  1457 => x"0c738f06",
  1458 => x"b7bc0ca0",
  1459 => x"5273bce0",
  1460 => x"082e0981",
  1461 => x"069838bc",
  1462 => x"dc08ff05",
  1463 => x"74327009",
  1464 => x"81057072",
  1465 => x"079f2a91",
  1466 => x"71315151",
  1467 => x"53537151",
  1468 => x"82ee2d81",
  1469 => x"14548e74",
  1470 => x"25c638b7",
  1471 => x"a8085271",
  1472 => x"b7ac0c02",
  1473 => x"94050d04",
  1474 => x"00ffffff",
  1475 => x"ff00ffff",
  1476 => x"ffff00ff",
  1477 => x"ffffff00",
  1478 => x"52657365",
  1479 => x"74000000",
  1480 => x"53617665",
  1481 => x"20616e64",
  1482 => x"20526573",
  1483 => x"65740000",
  1484 => x"4f707469",
  1485 => x"6f6e7320",
  1486 => x"10000000",
  1487 => x"536f756e",
  1488 => x"64201000",
  1489 => x"54757262",
  1490 => x"6f000000",
  1491 => x"4d6f7573",
  1492 => x"6520656d",
  1493 => x"756c6174",
  1494 => x"696f6e00",
  1495 => x"45786974",
  1496 => x"00000000",
  1497 => x"4d617374",
  1498 => x"65720000",
  1499 => x"4f504c4c",
  1500 => x"00000000",
  1501 => x"53434300",
  1502 => x"50534700",
  1503 => x"4261636b",
  1504 => x"00000000",
  1505 => x"5363616e",
  1506 => x"6c696e65",
  1507 => x"73000000",
  1508 => x"53442043",
  1509 => x"61726400",
  1510 => x"4a617061",
  1511 => x"6e657365",
  1512 => x"206b6579",
  1513 => x"206c6179",
  1514 => x"6f757400",
  1515 => x"32303438",
  1516 => x"4c422052",
  1517 => x"414d0000",
  1518 => x"34303936",
  1519 => x"4b422052",
  1520 => x"414d0000",
  1521 => x"536c323a",
  1522 => x"204e6f6e",
  1523 => x"65000000",
  1524 => x"536c323a",
  1525 => x"20455345",
  1526 => x"2d534343",
  1527 => x"20314d42",
  1528 => x"2f534343",
  1529 => x"2d490000",
  1530 => x"536c323a",
  1531 => x"20455345",
  1532 => x"2d52414d",
  1533 => x"20314d42",
  1534 => x"2f415343",
  1535 => x"49493800",
  1536 => x"536c323a",
  1537 => x"20455345",
  1538 => x"2d52414d",
  1539 => x"20314d42",
  1540 => x"2f415343",
  1541 => x"49493136",
  1542 => x"00000000",
  1543 => x"536c313a",
  1544 => x"204e6f6e",
  1545 => x"65000000",
  1546 => x"536c313a",
  1547 => x"20455345",
  1548 => x"2d534343",
  1549 => x"20314d42",
  1550 => x"2f534343",
  1551 => x"2d490000",
  1552 => x"536c313a",
  1553 => x"204d6567",
  1554 => x"6152414d",
  1555 => x"00000000",
  1556 => x"56474120",
  1557 => x"2d203331",
  1558 => x"4b487a2c",
  1559 => x"20363048",
  1560 => x"7a000000",
  1561 => x"56474120",
  1562 => x"2d203331",
  1563 => x"4b487a2c",
  1564 => x"20353048",
  1565 => x"7a000000",
  1566 => x"5456202d",
  1567 => x"20343830",
  1568 => x"692c2036",
  1569 => x"30487a00",
  1570 => x"496e6974",
  1571 => x"69616c69",
  1572 => x"7a696e67",
  1573 => x"20534420",
  1574 => x"63617264",
  1575 => x"0a000000",
  1576 => x"53444843",
  1577 => x"206e6f74",
  1578 => x"20737570",
  1579 => x"706f7274",
  1580 => x"65643b00",
  1581 => x"46617433",
  1582 => x"32206e6f",
  1583 => x"74207375",
  1584 => x"70706f72",
  1585 => x"7465643b",
  1586 => x"00000000",
  1587 => x"0a646973",
  1588 => x"61626c69",
  1589 => x"6e672053",
  1590 => x"44206361",
  1591 => x"72640a10",
  1592 => x"204f4b0a",
  1593 => x"00000000",
  1594 => x"4f434d53",
  1595 => x"58202020",
  1596 => x"43464700",
  1597 => x"54727969",
  1598 => x"6e67204d",
  1599 => x"53583342",
  1600 => x"494f532e",
  1601 => x"5359530a",
  1602 => x"00000000",
  1603 => x"4d535833",
  1604 => x"42494f53",
  1605 => x"53595300",
  1606 => x"54727969",
  1607 => x"6e672042",
  1608 => x"494f535f",
  1609 => x"4d32502e",
  1610 => x"524f4d0a",
  1611 => x"00000000",
  1612 => x"42494f53",
  1613 => x"5f4d3250",
  1614 => x"524f4d00",
  1615 => x"4c6f6164",
  1616 => x"696e6720",
  1617 => x"42494f53",
  1618 => x"0a000000",
  1619 => x"52656164",
  1620 => x"20666169",
  1621 => x"6c65640a",
  1622 => x"00000000",
  1623 => x"4c6f6164",
  1624 => x"696e6720",
  1625 => x"42494f53",
  1626 => x"20666169",
  1627 => x"6c65640a",
  1628 => x"00000000",
  1629 => x"4d425220",
  1630 => x"6661696c",
  1631 => x"0a000000",
  1632 => x"46415431",
  1633 => x"36202020",
  1634 => x"00000000",
  1635 => x"46415433",
  1636 => x"32202020",
  1637 => x"00000000",
  1638 => x"4e6f2070",
  1639 => x"61727469",
  1640 => x"74696f6e",
  1641 => x"20736967",
  1642 => x"0a000000",
  1643 => x"42616420",
  1644 => x"70617274",
  1645 => x"0a000000",
  1646 => x"53444843",
  1647 => x"20657272",
  1648 => x"6f72210a",
  1649 => x"00000000",
  1650 => x"53442069",
  1651 => x"6e69742e",
  1652 => x"2e2e0a00",
  1653 => x"53442063",
  1654 => x"61726420",
  1655 => x"72657365",
  1656 => x"74206661",
  1657 => x"696c6564",
  1658 => x"210a0000",
  1659 => x"57726974",
  1660 => x"65206661",
  1661 => x"696c6564",
  1662 => x"0a000000",
  1663 => x"16200000",
  1664 => x"14200000",
  1665 => x"15200000",
  1666 => x"00000002",
  1667 => x"00000002",
  1668 => x"00001718",
  1669 => x"00000666",
  1670 => x"00000002",
  1671 => x"00001720",
  1672 => x"00000658",
  1673 => x"00000004",
  1674 => x"00001730",
  1675 => x"00001ab4",
  1676 => x"00000004",
  1677 => x"0000173c",
  1678 => x"00001a6c",
  1679 => x"00000001",
  1680 => x"00001744",
  1681 => x"00000007",
  1682 => x"00000001",
  1683 => x"0000174c",
  1684 => x"0000000a",
  1685 => x"00000002",
  1686 => x"0000175c",
  1687 => x"000013c8",
  1688 => x"00000000",
  1689 => x"00000000",
  1690 => x"00000000",
  1691 => x"00000005",
  1692 => x"00001764",
  1693 => x"00000007",
  1694 => x"00000005",
  1695 => x"0000176c",
  1696 => x"00000007",
  1697 => x"00000005",
  1698 => x"00001774",
  1699 => x"00000007",
  1700 => x"00000005",
  1701 => x"00001778",
  1702 => x"00000007",
  1703 => x"00000004",
  1704 => x"0000177c",
  1705 => x"00001a0c",
  1706 => x"00000000",
  1707 => x"00000000",
  1708 => x"00000000",
  1709 => x"00000003",
  1710 => x"00001b44",
  1711 => x"00000003",
  1712 => x"00000001",
  1713 => x"00001784",
  1714 => x"0000000b",
  1715 => x"00000001",
  1716 => x"00001790",
  1717 => x"00000002",
  1718 => x"00000003",
  1719 => x"00001b38",
  1720 => x"00000003",
  1721 => x"00000003",
  1722 => x"00001b28",
  1723 => x"00000004",
  1724 => x"00000001",
  1725 => x"00001798",
  1726 => x"00000006",
  1727 => x"00000003",
  1728 => x"00001b20",
  1729 => x"00000002",
  1730 => x"00000004",
  1731 => x"0000177c",
  1732 => x"00001a0c",
  1733 => x"00000000",
  1734 => x"00000000",
  1735 => x"00000000",
  1736 => x"000017ac",
  1737 => x"000017b8",
  1738 => x"000017c4",
  1739 => x"000017d0",
  1740 => x"000017e8",
  1741 => x"00001800",
  1742 => x"0000181c",
  1743 => x"00001828",
  1744 => x"00001840",
  1745 => x"00001850",
  1746 => x"00001864",
  1747 => x"00001878",
  1748 => x"ffffffff",
  1749 => x"00000003",
  1750 => x"00000000",
  1751 => x"00000000",
  1752 => x"00000000",
  1753 => x"00000000",
  1754 => x"00000000",
  1755 => x"00000000",
  1756 => x"00000000",
  1757 => x"00000000",
  1758 => x"00000000",
  1759 => x"00000000",
  1760 => x"00000000",
  1761 => x"00000000",
  1762 => x"00000000",
  1763 => x"00000000",
  1764 => x"00000000",
  1765 => x"00000000",
  1766 => x"00000000",
  1767 => x"00000000",
  1768 => x"00000000",
  1769 => x"00000000",
  1770 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

