-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"000b0b0b",
     4 => x"0b8c04ff",
     5 => x"0d800404",
     6 => x"00000017",
     7 => x"00000000",
     8 => x"0b0b0bb7",
     9 => x"e8080b0b",
    10 => x"0bb7ec08",
    11 => x"0b0b0bb7",
    12 => x"f0080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"b7f00c0b",
    16 => x"0b0bb7ec",
    17 => x"0c0b0b0b",
    18 => x"b7e80c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0baec8",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"b7e870bd",
    57 => x"a0278b38",
    58 => x"80717084",
    59 => x"05530c81",
    60 => x"e2048c51",
    61 => x"8d8a0402",
    62 => x"fc050df8",
    63 => x"80518f0b",
    64 => x"b7f80c9f",
    65 => x"0bb7fc0c",
    66 => x"a0717081",
    67 => x"055334b7",
    68 => x"fc08ff05",
    69 => x"b7fc0cb7",
    70 => x"fc088025",
    71 => x"eb38b7f8",
    72 => x"08ff05b7",
    73 => x"f80cb7f8",
    74 => x"088025d7",
    75 => x"38028405",
    76 => x"0d0402f0",
    77 => x"050df880",
    78 => x"53f8a054",
    79 => x"83bf5273",
    80 => x"70810555",
    81 => x"33517073",
    82 => x"70810555",
    83 => x"34ff1252",
    84 => x"718025eb",
    85 => x"38fbc053",
    86 => x"9f52a073",
    87 => x"70810555",
    88 => x"34ff1252",
    89 => x"718025f2",
    90 => x"38029005",
    91 => x"0d0402f4",
    92 => x"050d7453",
    93 => x"8e0bb7f8",
    94 => x"08258f38",
    95 => x"82b22db7",
    96 => x"f808ff05",
    97 => x"b7f80c82",
    98 => x"f404b7f8",
    99 => x"08b7fc08",
   100 => x"5351728a",
   101 => x"2e098106",
   102 => x"b7387151",
   103 => x"719f24a0",
   104 => x"38b7f808",
   105 => x"a02911f8",
   106 => x"80115151",
   107 => x"a07134b7",
   108 => x"fc088105",
   109 => x"b7fc0cb7",
   110 => x"fc08519f",
   111 => x"7125e238",
   112 => x"800bb7fc",
   113 => x"0cb7f808",
   114 => x"8105b7f8",
   115 => x"0c83e404",
   116 => x"70a02912",
   117 => x"f8801151",
   118 => x"51727134",
   119 => x"b7fc0881",
   120 => x"05b7fc0c",
   121 => x"b7fc08a0",
   122 => x"2e098106",
   123 => x"8e38800b",
   124 => x"b7fc0cb7",
   125 => x"f8088105",
   126 => x"b7f80c02",
   127 => x"8c050d04",
   128 => x"02e8050d",
   129 => x"77795656",
   130 => x"880bfc16",
   131 => x"77712c8f",
   132 => x"06545254",
   133 => x"80537272",
   134 => x"25953871",
   135 => x"53fbe014",
   136 => x"51877134",
   137 => x"8114ff14",
   138 => x"545472f1",
   139 => x"387153f9",
   140 => x"1576712c",
   141 => x"87065351",
   142 => x"71802e8b",
   143 => x"38fbe014",
   144 => x"51717134",
   145 => x"81145472",
   146 => x"8e249538",
   147 => x"8f733153",
   148 => x"fbe01451",
   149 => x"a0713481",
   150 => x"14ff1454",
   151 => x"5472f138",
   152 => x"0298050d",
   153 => x"0402ec05",
   154 => x"0d800bb8",
   155 => x"800cf68c",
   156 => x"08f69008",
   157 => x"71882c56",
   158 => x"5481ff06",
   159 => x"52737225",
   160 => x"88387154",
   161 => x"820bb880",
   162 => x"0c72882c",
   163 => x"7381ff06",
   164 => x"54557473",
   165 => x"258b3872",
   166 => x"b8800884",
   167 => x"07b8800c",
   168 => x"5573842b",
   169 => x"86a07125",
   170 => x"83713170",
   171 => x"0b0b0bb4",
   172 => x"c80c8171",
   173 => x"2bff05f6",
   174 => x"880cfecc",
   175 => x"13ff122c",
   176 => x"788829ff",
   177 => x"94057081",
   178 => x"2cb88008",
   179 => x"52585255",
   180 => x"51525476",
   181 => x"802e8538",
   182 => x"70810751",
   183 => x"70f6940c",
   184 => x"71098105",
   185 => x"f6800c72",
   186 => x"098105f6",
   187 => x"840c0294",
   188 => x"050d0402",
   189 => x"f4050d74",
   190 => x"53727081",
   191 => x"055480f5",
   192 => x"2d527180",
   193 => x"2e893871",
   194 => x"5182ee2d",
   195 => x"85f90402",
   196 => x"8c050d04",
   197 => x"02f8050d",
   198 => x"a5ff2d80",
   199 => x"da51a7b6",
   200 => x"2db7e808",
   201 => x"812a7081",
   202 => x"06515271",
   203 => x"802ee938",
   204 => x"0288050d",
   205 => x"0402f405",
   206 => x"0dbd9008",
   207 => x"99c406b6",
   208 => x"c40b80f5",
   209 => x"2d525270",
   210 => x"802e8638",
   211 => x"71848007",
   212 => x"52b5fc0b",
   213 => x"80f52d72",
   214 => x"07b6a00b",
   215 => x"80f52d70",
   216 => x"812a7081",
   217 => x"06515354",
   218 => x"5270802e",
   219 => x"86387182",
   220 => x"80075272",
   221 => x"81065170",
   222 => x"802e8538",
   223 => x"71880752",
   224 => x"b6ac0b80",
   225 => x"f52d7084",
   226 => x"2b730781",
   227 => x"8432b7e8",
   228 => x"0c51028c",
   229 => x"050d0402",
   230 => x"f4050d74",
   231 => x"70818432",
   232 => x"bd900c70",
   233 => x"83065253",
   234 => x"70b5f40b",
   235 => x"880581b7",
   236 => x"2d72892a",
   237 => x"70810651",
   238 => x"5170b6c4",
   239 => x"0b81b72d",
   240 => x"72832a81",
   241 => x"0673882a",
   242 => x"70810651",
   243 => x"52527080",
   244 => x"2e853871",
   245 => x"82075271",
   246 => x"b6a00b81",
   247 => x"b72d7284",
   248 => x"2c708306",
   249 => x"515170b6",
   250 => x"ac0b81b7",
   251 => x"2d70b7e8",
   252 => x"0c028c05",
   253 => x"0d0402f4",
   254 => x"050db5ac",
   255 => x"0b881180",
   256 => x"f52d8c12",
   257 => x"881180f5",
   258 => x"2d70842b",
   259 => x"73078c13",
   260 => x"881180f5",
   261 => x"2d70882b",
   262 => x"73079413",
   263 => x"80f52d70",
   264 => x"8c2b7207",
   265 => x"b7e80c53",
   266 => x"53535353",
   267 => x"56525351",
   268 => x"028c050d",
   269 => x"0402f405",
   270 => x"0d74b5ac",
   271 => x"71870655",
   272 => x"53517288",
   273 => x"1381b72d",
   274 => x"8c127184",
   275 => x"2c708706",
   276 => x"55525272",
   277 => x"881381b7",
   278 => x"2d8c1271",
   279 => x"842c7087",
   280 => x"06555252",
   281 => x"72881381",
   282 => x"b72d7084",
   283 => x"2c708706",
   284 => x"51517094",
   285 => x"1381b72d",
   286 => x"028c050d",
   287 => x"0402d405",
   288 => x"0d7cb1c8",
   289 => x"525585f3",
   290 => x"2d9db02d",
   291 => x"b7e80880",
   292 => x"2e839d38",
   293 => x"86b52db7",
   294 => x"e808538f",
   295 => x"f92db7e8",
   296 => x"0854b7e8",
   297 => x"08802e83",
   298 => x"8938a1b3",
   299 => x"2db7e808",
   300 => x"802e8738",
   301 => x"b1e05189",
   302 => x"c704999c",
   303 => x"2db7e808",
   304 => x"802ea238",
   305 => x"b1f45185",
   306 => x"f32db28c",
   307 => x"5185f32d",
   308 => x"86942d72",
   309 => x"84075381",
   310 => x"0bfec40c",
   311 => x"72fec00c",
   312 => x"72518797",
   313 => x"2d840bfe",
   314 => x"c40cb2a8",
   315 => x"52b88851",
   316 => x"968b2db7",
   317 => x"e808802e",
   318 => x"80dc3874",
   319 => x"822e0981",
   320 => x"06af3872",
   321 => x"b8940c87",
   322 => x"f62db7e8",
   323 => x"08b8980c",
   324 => x"b89c5480",
   325 => x"fd538074",
   326 => x"70840556",
   327 => x"0cff1353",
   328 => x"728025f2",
   329 => x"38b89452",
   330 => x"b8885198",
   331 => x"f62d8ad6",
   332 => x"0474812e",
   333 => x"0981069e",
   334 => x"38b89452",
   335 => x"b8885198",
   336 => x"d02db894",
   337 => x"08b89808",
   338 => x"525388b5",
   339 => x"2d72fec0",
   340 => x"0c725187",
   341 => x"972db2b4",
   342 => x"5185f32d",
   343 => x"b2cc52b8",
   344 => x"8851968b",
   345 => x"2db7e808",
   346 => x"9838b2d8",
   347 => x"5185f32d",
   348 => x"b2f052b8",
   349 => x"8851968b",
   350 => x"2db7e808",
   351 => x"802e81b0",
   352 => x"38b2fc51",
   353 => x"85f32db8",
   354 => x"8c085780",
   355 => x"77595a76",
   356 => x"7a2e8b38",
   357 => x"811a7881",
   358 => x"2a595a77",
   359 => x"f738f71a",
   360 => x"5a807725",
   361 => x"81803879",
   362 => x"52775184",
   363 => x"802db894",
   364 => x"52b88851",
   365 => x"98d02db7",
   366 => x"e80853b7",
   367 => x"e808802e",
   368 => x"80c938b8",
   369 => x"945b8059",
   370 => x"8bf8047a",
   371 => x"7084055c",
   372 => x"087081ff",
   373 => x"0671882c",
   374 => x"7081ff06",
   375 => x"73902c70",
   376 => x"81ff0675",
   377 => x"982afec8",
   378 => x"0cfec80c",
   379 => x"58fec80c",
   380 => x"57fec80c",
   381 => x"841a5a53",
   382 => x"76538480",
   383 => x"77258438",
   384 => x"84805372",
   385 => x"7924c438",
   386 => x"8c9604b3",
   387 => x"8c5185f3",
   388 => x"2d72548c",
   389 => x"b204b888",
   390 => x"5198a32d",
   391 => x"fc801781",
   392 => x"1959578b",
   393 => x"a104820b",
   394 => x"fec40c81",
   395 => x"548cb204",
   396 => x"805473b7",
   397 => x"e80c02ac",
   398 => x"050d0402",
   399 => x"f8050da8",
   400 => x"862d81f7",
   401 => x"2d815184",
   402 => x"e52dfec4",
   403 => x"5281720c",
   404 => x"a4ff2da4",
   405 => x"ff2d8472",
   406 => x"0c735188",
   407 => x"fd2db4cc",
   408 => x"51a9e42d",
   409 => x"805184e5",
   410 => x"2d028805",
   411 => x"0d0402fc",
   412 => x"050d8251",
   413 => x"8cbb2d02",
   414 => x"84050d04",
   415 => x"02fc050d",
   416 => x"80518cbb",
   417 => x"2d028405",
   418 => x"0d0402ec",
   419 => x"050d84b8",
   420 => x"5187972d",
   421 => x"810bfec4",
   422 => x"0c84b80b",
   423 => x"fec00c84",
   424 => x"0bfec40c",
   425 => x"830bfecc",
   426 => x"0ca59a2d",
   427 => x"a7fa2da4",
   428 => x"ff2da4ff",
   429 => x"2d81f72d",
   430 => x"815184e5",
   431 => x"2da4ff2d",
   432 => x"a4ff2d81",
   433 => x"5184e52d",
   434 => x"815188fd",
   435 => x"2db7e808",
   436 => x"802e81d2",
   437 => x"38805184",
   438 => x"e52db4cc",
   439 => x"51a9e42d",
   440 => x"bcf00889",
   441 => x"38bcf408",
   442 => x"802e80e2",
   443 => x"38fed008",
   444 => x"70810651",
   445 => x"5271802e",
   446 => x"80d438a8",
   447 => x"802dbcf0",
   448 => x"0870bcf4",
   449 => x"08705755",
   450 => x"565280ff",
   451 => x"72258438",
   452 => x"80ff5280",
   453 => x"ff732584",
   454 => x"3880ff53",
   455 => x"71ff8025",
   456 => x"8438ff80",
   457 => x"5272ff80",
   458 => x"258438ff",
   459 => x"80537472",
   460 => x"31bcf00c",
   461 => x"737331bc",
   462 => x"f40ca7fa",
   463 => x"2d71882b",
   464 => x"83fe8006",
   465 => x"7381ff06",
   466 => x"7107fed0",
   467 => x"0c52a5ff",
   468 => x"2da9f42d",
   469 => x"b7e80853",
   470 => x"86b52db7",
   471 => x"e808fec0",
   472 => x"0c87f62d",
   473 => x"b7e808fe",
   474 => x"d40c86b5",
   475 => x"2db7e808",
   476 => x"b884082e",
   477 => x"9c38b7e8",
   478 => x"08b8840c",
   479 => x"84527251",
   480 => x"84e52da4",
   481 => x"ff2da4ff",
   482 => x"2dff1252",
   483 => x"718025ee",
   484 => x"3872802e",
   485 => x"89388a0b",
   486 => x"fec40c8d",
   487 => x"e004820b",
   488 => x"fec40c8d",
   489 => x"e004b39c",
   490 => x"5185f32d",
   491 => x"820bfec4",
   492 => x"0c800bb7",
   493 => x"e80c0294",
   494 => x"050d0402",
   495 => x"e8050d77",
   496 => x"797b5855",
   497 => x"55805372",
   498 => x"7625a338",
   499 => x"74708105",
   500 => x"5680f52d",
   501 => x"74708105",
   502 => x"5680f52d",
   503 => x"52527171",
   504 => x"2e863881",
   505 => x"518ff004",
   506 => x"8113538f",
   507 => x"c7048051",
   508 => x"70b7e80c",
   509 => x"0298050d",
   510 => x"0402d805",
   511 => x"0d800bbc",
   512 => x"9c0cb894",
   513 => x"528051a0",
   514 => x"982db7e8",
   515 => x"0854b7e8",
   516 => x"088c38b3",
   517 => x"b45185f3",
   518 => x"2d735595",
   519 => x"94048056",
   520 => x"810bbcc0",
   521 => x"0c8853b3",
   522 => x"c052b8ca",
   523 => x"518fbb2d",
   524 => x"b7e80876",
   525 => x"2e098106",
   526 => x"8738b7e8",
   527 => x"08bcc00c",
   528 => x"8853b3cc",
   529 => x"52b8e651",
   530 => x"8fbb2db7",
   531 => x"e8088738",
   532 => x"b7e808bc",
   533 => x"c00cbcc0",
   534 => x"08802e80",
   535 => x"f638bbda",
   536 => x"0b80f52d",
   537 => x"bbdb0b80",
   538 => x"f52d7198",
   539 => x"2b71902b",
   540 => x"07bbdc0b",
   541 => x"80f52d70",
   542 => x"882b7207",
   543 => x"bbdd0b80",
   544 => x"f52d7107",
   545 => x"bc920b80",
   546 => x"f52dbc93",
   547 => x"0b80f52d",
   548 => x"71882b07",
   549 => x"535f5452",
   550 => x"5a565755",
   551 => x"7381abaa",
   552 => x"2e098106",
   553 => x"8d387551",
   554 => x"a1ba2db7",
   555 => x"e8085691",
   556 => x"bf047382",
   557 => x"d4d52e87",
   558 => x"38b3d851",
   559 => x"928004b8",
   560 => x"94527551",
   561 => x"a0982db7",
   562 => x"e80855b7",
   563 => x"e808802e",
   564 => x"83c23888",
   565 => x"53b3cc52",
   566 => x"b8e6518f",
   567 => x"bb2db7e8",
   568 => x"08893881",
   569 => x"0bbc9c0c",
   570 => x"92860488",
   571 => x"53b3c052",
   572 => x"b8ca518f",
   573 => x"bb2db7e8",
   574 => x"08802e8a",
   575 => x"38b3ec51",
   576 => x"85f32d92",
   577 => x"e004bc92",
   578 => x"0b80f52d",
   579 => x"547380d5",
   580 => x"2e098106",
   581 => x"80ca38bc",
   582 => x"930b80f5",
   583 => x"2d547381",
   584 => x"aa2e0981",
   585 => x"06ba3880",
   586 => x"0bb8940b",
   587 => x"80f52d56",
   588 => x"547481e9",
   589 => x"2e833881",
   590 => x"547481eb",
   591 => x"2e8c3880",
   592 => x"5573752e",
   593 => x"09810682",
   594 => x"cb38b89f",
   595 => x"0b80f52d",
   596 => x"55748d38",
   597 => x"b8a00b80",
   598 => x"f52d5473",
   599 => x"822e8638",
   600 => x"80559594",
   601 => x"04b8a10b",
   602 => x"80f52d70",
   603 => x"bc940cff",
   604 => x"05bc980c",
   605 => x"b8a20b80",
   606 => x"f52db8a3",
   607 => x"0b80f52d",
   608 => x"58760577",
   609 => x"82802905",
   610 => x"70bca00c",
   611 => x"b8a40b80",
   612 => x"f52d70bc",
   613 => x"b40cbc9c",
   614 => x"08595758",
   615 => x"76802e81",
   616 => x"a3388853",
   617 => x"b3cc52b8",
   618 => x"e6518fbb",
   619 => x"2db7e808",
   620 => x"81e238bc",
   621 => x"94087084",
   622 => x"2bbcb80c",
   623 => x"70bcb00c",
   624 => x"b8b90b80",
   625 => x"f52db8b8",
   626 => x"0b80f52d",
   627 => x"71828029",
   628 => x"05b8ba0b",
   629 => x"80f52d70",
   630 => x"84808029",
   631 => x"12b8bb0b",
   632 => x"80f52d70",
   633 => x"81800a29",
   634 => x"1270bcbc",
   635 => x"0cbcb408",
   636 => x"7129bca0",
   637 => x"080570bc",
   638 => x"a40cb8c1",
   639 => x"0b80f52d",
   640 => x"b8c00b80",
   641 => x"f52d7182",
   642 => x"802905b8",
   643 => x"c20b80f5",
   644 => x"2d708480",
   645 => x"802912b8",
   646 => x"c30b80f5",
   647 => x"2d70982b",
   648 => x"81f00a06",
   649 => x"720570bc",
   650 => x"a80cfe11",
   651 => x"7e297705",
   652 => x"bcac0c52",
   653 => x"59524354",
   654 => x"5e515259",
   655 => x"525d5759",
   656 => x"57959204",
   657 => x"b8a60b80",
   658 => x"f52db8a5",
   659 => x"0b80f52d",
   660 => x"71828029",
   661 => x"0570bcb8",
   662 => x"0c70a029",
   663 => x"83ff0570",
   664 => x"892a70bc",
   665 => x"b00cb8ab",
   666 => x"0b80f52d",
   667 => x"b8aa0b80",
   668 => x"f52d7182",
   669 => x"80290570",
   670 => x"bcbc0c7b",
   671 => x"71291e70",
   672 => x"bcac0c7d",
   673 => x"bca80c73",
   674 => x"05bca40c",
   675 => x"555e5151",
   676 => x"55558155",
   677 => x"74b7e80c",
   678 => x"02a8050d",
   679 => x"0402ec05",
   680 => x"0d767087",
   681 => x"2c7180ff",
   682 => x"06555654",
   683 => x"bc9c088a",
   684 => x"3873882c",
   685 => x"7481ff06",
   686 => x"5455b894",
   687 => x"52bca008",
   688 => x"1551a098",
   689 => x"2db7e808",
   690 => x"54b7e808",
   691 => x"802eb338",
   692 => x"bc9c0880",
   693 => x"2e983872",
   694 => x"8429b894",
   695 => x"05700852",
   696 => x"53a1ba2d",
   697 => x"b7e808f0",
   698 => x"0a065396",
   699 => x"80047210",
   700 => x"b8940570",
   701 => x"80e02d52",
   702 => x"53a1ea2d",
   703 => x"b7e80853",
   704 => x"725473b7",
   705 => x"e80c0294",
   706 => x"050d0402",
   707 => x"c8050d7f",
   708 => x"615f5b80",
   709 => x"0bbca808",
   710 => x"bcac0859",
   711 => x"5d56bc9c",
   712 => x"08762e8a",
   713 => x"38bc9408",
   714 => x"842b5896",
   715 => x"b404bcb0",
   716 => x"08842b58",
   717 => x"80597878",
   718 => x"2781a938",
   719 => x"788f06a0",
   720 => x"17575473",
   721 => x"8f38b894",
   722 => x"52765181",
   723 => x"1757a098",
   724 => x"2db89456",
   725 => x"807680f5",
   726 => x"2d565474",
   727 => x"742e8338",
   728 => x"81547481",
   729 => x"e52e80f6",
   730 => x"38817075",
   731 => x"06555d73",
   732 => x"802e80ea",
   733 => x"388b1680",
   734 => x"f52d9806",
   735 => x"5a7980de",
   736 => x"388b537d",
   737 => x"5275518f",
   738 => x"bb2db7e8",
   739 => x"0880cf38",
   740 => x"9c160851",
   741 => x"a1ba2db7",
   742 => x"e808841c",
   743 => x"0c9a1680",
   744 => x"e02d51a1",
   745 => x"ea2db7e8",
   746 => x"08b7e808",
   747 => x"881d0cb7",
   748 => x"e8085555",
   749 => x"bc9c0880",
   750 => x"2e983894",
   751 => x"1680e02d",
   752 => x"51a1ea2d",
   753 => x"b7e80890",
   754 => x"2b83fff0",
   755 => x"0a067016",
   756 => x"51547388",
   757 => x"1c0c797b",
   758 => x"0c7c5498",
   759 => x"9a048119",
   760 => x"5996b604",
   761 => x"bc9c0880",
   762 => x"2eae387b",
   763 => x"51959d2d",
   764 => x"b7e808b7",
   765 => x"e80880ff",
   766 => x"fffff806",
   767 => x"555c7380",
   768 => x"fffffff8",
   769 => x"2e9238b7",
   770 => x"e808fe05",
   771 => x"bc940829",
   772 => x"bca40805",
   773 => x"5796b404",
   774 => x"805473b7",
   775 => x"e80c02b8",
   776 => x"050d0402",
   777 => x"f4050d74",
   778 => x"70088105",
   779 => x"710c7008",
   780 => x"bc980806",
   781 => x"5353718e",
   782 => x"38881308",
   783 => x"51959d2d",
   784 => x"b7e80888",
   785 => x"140c810b",
   786 => x"b7e80c02",
   787 => x"8c050d04",
   788 => x"02f0050d",
   789 => x"75881108",
   790 => x"fe05bc94",
   791 => x"0829bca4",
   792 => x"08117208",
   793 => x"bc980806",
   794 => x"05795553",
   795 => x"5454a098",
   796 => x"2d029005",
   797 => x"0d0402f0",
   798 => x"050d7588",
   799 => x"1108fe05",
   800 => x"bc940829",
   801 => x"bca40811",
   802 => x"7208bc98",
   803 => x"08060579",
   804 => x"55535454",
   805 => x"9ed82d02",
   806 => x"90050d04",
   807 => x"bc9c08b7",
   808 => x"e80c0402",
   809 => x"f4050dd4",
   810 => x"5281ff72",
   811 => x"0c710853",
   812 => x"81ff720c",
   813 => x"72882b83",
   814 => x"fe800672",
   815 => x"087081ff",
   816 => x"06515253",
   817 => x"81ff720c",
   818 => x"72710788",
   819 => x"2b720870",
   820 => x"81ff0651",
   821 => x"525381ff",
   822 => x"720c7271",
   823 => x"07882b72",
   824 => x"087081ff",
   825 => x"067207b7",
   826 => x"e80c5253",
   827 => x"028c050d",
   828 => x"0402f405",
   829 => x"0d747671",
   830 => x"81ff06d4",
   831 => x"0c5353bc",
   832 => x"c4088538",
   833 => x"71892b52",
   834 => x"71982ad4",
   835 => x"0c71902a",
   836 => x"7081ff06",
   837 => x"d40c5171",
   838 => x"882a7081",
   839 => x"ff06d40c",
   840 => x"517181ff",
   841 => x"06d40c72",
   842 => x"902a7081",
   843 => x"ff06d40c",
   844 => x"51d40870",
   845 => x"81ff0651",
   846 => x"5182b8bf",
   847 => x"527081ff",
   848 => x"2e098106",
   849 => x"943881ff",
   850 => x"0bd40cd4",
   851 => x"087081ff",
   852 => x"06ff1454",
   853 => x"515171e5",
   854 => x"3870b7e8",
   855 => x"0c028c05",
   856 => x"0d0402fc",
   857 => x"050d81c7",
   858 => x"5181ff0b",
   859 => x"d40cff11",
   860 => x"51708025",
   861 => x"f4380284",
   862 => x"050d0402",
   863 => x"f0050d9a",
   864 => x"e22d8fcf",
   865 => x"53805287",
   866 => x"fc80f751",
   867 => x"99f12db7",
   868 => x"e80854b7",
   869 => x"e808812e",
   870 => x"098106a3",
   871 => x"3881ff0b",
   872 => x"d40c820a",
   873 => x"52849c80",
   874 => x"e95199f1",
   875 => x"2db7e808",
   876 => x"8b3881ff",
   877 => x"0bd40c73",
   878 => x"539bc504",
   879 => x"9ae22dff",
   880 => x"135372c1",
   881 => x"3872b7e8",
   882 => x"0c029005",
   883 => x"0d0402f4",
   884 => x"050d81ff",
   885 => x"0bd40c93",
   886 => x"53805287",
   887 => x"fc80c151",
   888 => x"99f12db7",
   889 => x"e8088b38",
   890 => x"81ff0bd4",
   891 => x"0c81539b",
   892 => x"fb049ae2",
   893 => x"2dff1353",
   894 => x"72df3872",
   895 => x"b7e80c02",
   896 => x"8c050d04",
   897 => x"02f0050d",
   898 => x"9ae22d83",
   899 => x"aa52849c",
   900 => x"80c85199",
   901 => x"f12db7e8",
   902 => x"08812e09",
   903 => x"81069238",
   904 => x"99a32db7",
   905 => x"e80883ff",
   906 => x"ff065372",
   907 => x"83aa2e97",
   908 => x"389bce2d",
   909 => x"9cc20481",
   910 => x"549da704",
   911 => x"b3f85185",
   912 => x"f32d8054",
   913 => x"9da70481",
   914 => x"ff0bd40c",
   915 => x"b1539afb",
   916 => x"2db7e808",
   917 => x"802e80c0",
   918 => x"38805287",
   919 => x"fc80fa51",
   920 => x"99f12db7",
   921 => x"e808b138",
   922 => x"81ff0bd4",
   923 => x"0cd40853",
   924 => x"81ff0bd4",
   925 => x"0c81ff0b",
   926 => x"d40c81ff",
   927 => x"0bd40c81",
   928 => x"ff0bd40c",
   929 => x"72862a70",
   930 => x"8106b7e8",
   931 => x"08565153",
   932 => x"72802e93",
   933 => x"389cb704",
   934 => x"72822eff",
   935 => x"9f38ff13",
   936 => x"5372ffaa",
   937 => x"38725473",
   938 => x"b7e80c02",
   939 => x"90050d04",
   940 => x"02f0050d",
   941 => x"810bbcc4",
   942 => x"0c8454d0",
   943 => x"08708f2a",
   944 => x"70810651",
   945 => x"515372f3",
   946 => x"3872d00c",
   947 => x"9ae22db4",
   948 => x"885185f3",
   949 => x"2dd00870",
   950 => x"8f2a7081",
   951 => x"06515153",
   952 => x"72f33881",
   953 => x"0bd00cb1",
   954 => x"53805284",
   955 => x"d480c051",
   956 => x"99f12db7",
   957 => x"e808812e",
   958 => x"a1387282",
   959 => x"2e098106",
   960 => x"8c38b494",
   961 => x"5185f32d",
   962 => x"80539ecf",
   963 => x"04ff1353",
   964 => x"72d738ff",
   965 => x"145473ff",
   966 => x"a2389c84",
   967 => x"2db7e808",
   968 => x"bcc40cb7",
   969 => x"e8088b38",
   970 => x"815287fc",
   971 => x"80d05199",
   972 => x"f12d81ff",
   973 => x"0bd40cd0",
   974 => x"08708f2a",
   975 => x"70810651",
   976 => x"515372f3",
   977 => x"3872d00c",
   978 => x"81ff0bd4",
   979 => x"0c815372",
   980 => x"b7e80c02",
   981 => x"90050d04",
   982 => x"02e8050d",
   983 => x"785681ff",
   984 => x"0bd40cd0",
   985 => x"08708f2a",
   986 => x"70810651",
   987 => x"515372f3",
   988 => x"3882810b",
   989 => x"d00c81ff",
   990 => x"0bd40c77",
   991 => x"5287fc80",
   992 => x"d85199f1",
   993 => x"2db7e808",
   994 => x"802e8c38",
   995 => x"b4ac5185",
   996 => x"f32d8153",
   997 => x"a08f0481",
   998 => x"ff0bd40c",
   999 => x"81fe0bd4",
  1000 => x"0c80ff55",
  1001 => x"75708405",
  1002 => x"57087098",
  1003 => x"2ad40c70",
  1004 => x"902c7081",
  1005 => x"ff06d40c",
  1006 => x"5470882c",
  1007 => x"7081ff06",
  1008 => x"d40c5470",
  1009 => x"81ff06d4",
  1010 => x"0c54ff15",
  1011 => x"55748025",
  1012 => x"d33881ff",
  1013 => x"0bd40c81",
  1014 => x"ff0bd40c",
  1015 => x"81ff0bd4",
  1016 => x"0c868da0",
  1017 => x"5481ff0b",
  1018 => x"d40cd408",
  1019 => x"81ff0655",
  1020 => x"748738ff",
  1021 => x"145473ed",
  1022 => x"3881ff0b",
  1023 => x"d40cd008",
  1024 => x"708f2a70",
  1025 => x"81065151",
  1026 => x"5372f338",
  1027 => x"72d00c72",
  1028 => x"b7e80c02",
  1029 => x"98050d04",
  1030 => x"02e8050d",
  1031 => x"78558056",
  1032 => x"81ff0bd4",
  1033 => x"0cd00870",
  1034 => x"8f2a7081",
  1035 => x"06515153",
  1036 => x"72f33882",
  1037 => x"810bd00c",
  1038 => x"81ff0bd4",
  1039 => x"0c775287",
  1040 => x"fc80d151",
  1041 => x"99f12d80",
  1042 => x"dbc6df54",
  1043 => x"b7e80880",
  1044 => x"2e8a38b3",
  1045 => x"8c5185f3",
  1046 => x"2da1aa04",
  1047 => x"81ff0bd4",
  1048 => x"0cd40870",
  1049 => x"81ff0651",
  1050 => x"537281fe",
  1051 => x"2e098106",
  1052 => x"9d3880ff",
  1053 => x"5399a32d",
  1054 => x"b7e80875",
  1055 => x"70840557",
  1056 => x"0cff1353",
  1057 => x"728025ed",
  1058 => x"388156a1",
  1059 => x"9404ff14",
  1060 => x"5473c938",
  1061 => x"81ff0bd4",
  1062 => x"0cd00870",
  1063 => x"8f2a7081",
  1064 => x"06515153",
  1065 => x"72f33872",
  1066 => x"d00c75b7",
  1067 => x"e80c0298",
  1068 => x"050d04bc",
  1069 => x"c408b7e8",
  1070 => x"0c0402f4",
  1071 => x"050d7470",
  1072 => x"882a83fe",
  1073 => x"80067072",
  1074 => x"982a0772",
  1075 => x"882b87fc",
  1076 => x"80800673",
  1077 => x"982b81f0",
  1078 => x"0a067173",
  1079 => x"0707b7e8",
  1080 => x"0c565153",
  1081 => x"51028c05",
  1082 => x"0d0402f8",
  1083 => x"050d028e",
  1084 => x"0580f52d",
  1085 => x"74882b07",
  1086 => x"7083ffff",
  1087 => x"06b7e80c",
  1088 => x"51028805",
  1089 => x"0d0402fc",
  1090 => x"050d7251",
  1091 => x"80710c80",
  1092 => x"0b84120c",
  1093 => x"0284050d",
  1094 => x"0402f005",
  1095 => x"0d757008",
  1096 => x"84120853",
  1097 => x"5353ff54",
  1098 => x"71712ea8",
  1099 => x"38a8802d",
  1100 => x"84130870",
  1101 => x"84291488",
  1102 => x"11700870",
  1103 => x"81ff0684",
  1104 => x"18088111",
  1105 => x"8706841a",
  1106 => x"0c535155",
  1107 => x"515151a7",
  1108 => x"fa2d7154",
  1109 => x"73b7e80c",
  1110 => x"0290050d",
  1111 => x"0402f405",
  1112 => x"0da8802d",
  1113 => x"e008e408",
  1114 => x"718b2a70",
  1115 => x"81065153",
  1116 => x"54527080",
  1117 => x"2e9d38bc",
  1118 => x"c8087084",
  1119 => x"29bcd005",
  1120 => x"7381ff06",
  1121 => x"710c5151",
  1122 => x"bcc80881",
  1123 => x"118706bc",
  1124 => x"c80c5172",
  1125 => x"8b2a7081",
  1126 => x"06515170",
  1127 => x"802e8192",
  1128 => x"38b79808",
  1129 => x"8429bcfc",
  1130 => x"057381ff",
  1131 => x"06710c51",
  1132 => x"b7980881",
  1133 => x"05b7980c",
  1134 => x"850bb794",
  1135 => x"0cb79808",
  1136 => x"b790082e",
  1137 => x"09810681",
  1138 => x"a638800b",
  1139 => x"b7980cbd",
  1140 => x"8c08819b",
  1141 => x"38bcfc08",
  1142 => x"70097083",
  1143 => x"06fecc0c",
  1144 => x"5270852a",
  1145 => x"708106bc",
  1146 => x"f4085551",
  1147 => x"52537080",
  1148 => x"2e8e38bd",
  1149 => x"8408fe80",
  1150 => x"3212bcf4",
  1151 => x"0ca48704",
  1152 => x"bd840812",
  1153 => x"bcf40c72",
  1154 => x"842a7081",
  1155 => x"06bcf008",
  1156 => x"54515170",
  1157 => x"802e9038",
  1158 => x"bd800881",
  1159 => x"ff321281",
  1160 => x"05bcf00c",
  1161 => x"a4ef0471",
  1162 => x"bd800831",
  1163 => x"bcf00ca4",
  1164 => x"ef04b794",
  1165 => x"08ff05b7",
  1166 => x"940cb794",
  1167 => x"08ff2e09",
  1168 => x"8106ac38",
  1169 => x"b7980880",
  1170 => x"2e923881",
  1171 => x"0bbd8c0c",
  1172 => x"870bb790",
  1173 => x"0831b790",
  1174 => x"0ca4ea04",
  1175 => x"bd8c0851",
  1176 => x"70802e86",
  1177 => x"38ff11bd",
  1178 => x"8c0c800b",
  1179 => x"b7980c80",
  1180 => x"0bbcf80c",
  1181 => x"a7f32da7",
  1182 => x"fa2d028c",
  1183 => x"050d0402",
  1184 => x"fc050da8",
  1185 => x"802d810b",
  1186 => x"bcf80ca7",
  1187 => x"fa2dbcf8",
  1188 => x"085170fa",
  1189 => x"38028405",
  1190 => x"0d0402f8",
  1191 => x"050dbcc8",
  1192 => x"51a2862d",
  1193 => x"800bbd8c",
  1194 => x"0c830bb7",
  1195 => x"900ce408",
  1196 => x"708c2a70",
  1197 => x"81065151",
  1198 => x"5271802e",
  1199 => x"8638840b",
  1200 => x"b7900ce4",
  1201 => x"08708d2a",
  1202 => x"70810651",
  1203 => x"51527180",
  1204 => x"2e9f3887",
  1205 => x"0bb79008",
  1206 => x"31b7900c",
  1207 => x"e408708a",
  1208 => x"2a708106",
  1209 => x"51515271",
  1210 => x"802ef138",
  1211 => x"81f40be4",
  1212 => x"0ca2dd51",
  1213 => x"a7ef2da7",
  1214 => x"992d0288",
  1215 => x"050d0402",
  1216 => x"f4050da7",
  1217 => x"8104b7e8",
  1218 => x"0881f02e",
  1219 => x"09810689",
  1220 => x"38810bb7",
  1221 => x"dc0ca781",
  1222 => x"04b7e808",
  1223 => x"81e02e09",
  1224 => x"81068938",
  1225 => x"810bb7e0",
  1226 => x"0ca78104",
  1227 => x"b7e80852",
  1228 => x"b7e00880",
  1229 => x"2e8838b7",
  1230 => x"e8088180",
  1231 => x"05527184",
  1232 => x"2c728f06",
  1233 => x"5353b7dc",
  1234 => x"08802e99",
  1235 => x"38728429",
  1236 => x"b79c0572",
  1237 => x"1381712b",
  1238 => x"70097308",
  1239 => x"06730c51",
  1240 => x"5353a6f7",
  1241 => x"04728429",
  1242 => x"b79c0572",
  1243 => x"1383712b",
  1244 => x"72080772",
  1245 => x"0c535380",
  1246 => x"0bb7e00c",
  1247 => x"800bb7dc",
  1248 => x"0cbcc851",
  1249 => x"a2992db7",
  1250 => x"e808ff24",
  1251 => x"fef83880",
  1252 => x"0bb7e80c",
  1253 => x"028c050d",
  1254 => x"0402f805",
  1255 => x"0db79c52",
  1256 => x"8f518072",
  1257 => x"70840554",
  1258 => x"0cff1151",
  1259 => x"708025f2",
  1260 => x"38028805",
  1261 => x"0d0402f0",
  1262 => x"050d7551",
  1263 => x"a8802d70",
  1264 => x"822cfc06",
  1265 => x"b79c1172",
  1266 => x"109e0671",
  1267 => x"0870722a",
  1268 => x"70830682",
  1269 => x"742b7009",
  1270 => x"7406760c",
  1271 => x"54515657",
  1272 => x"535153a7",
  1273 => x"fa2d71b7",
  1274 => x"e80c0290",
  1275 => x"050d0471",
  1276 => x"980c04ff",
  1277 => x"b008b7e8",
  1278 => x"0c04810b",
  1279 => x"ffb00c04",
  1280 => x"800bffb0",
  1281 => x"0c0402fc",
  1282 => x"050d800b",
  1283 => x"b7e40c80",
  1284 => x"5184e52d",
  1285 => x"0284050d",
  1286 => x"0402ec05",
  1287 => x"0d765480",
  1288 => x"52870b88",
  1289 => x"1580f52d",
  1290 => x"56537472",
  1291 => x"248338a0",
  1292 => x"53725182",
  1293 => x"ee2d8112",
  1294 => x"8b1580f5",
  1295 => x"2d545272",
  1296 => x"7225de38",
  1297 => x"0294050d",
  1298 => x"0402f005",
  1299 => x"0dbd9408",
  1300 => x"5481f72d",
  1301 => x"800bbd98",
  1302 => x"0c730880",
  1303 => x"2e818038",
  1304 => x"820bb7fc",
  1305 => x"0cbd9808",
  1306 => x"8f06b7f8",
  1307 => x"0c730852",
  1308 => x"71832e96",
  1309 => x"38718326",
  1310 => x"89387181",
  1311 => x"2eaf38a9",
  1312 => x"ca047185",
  1313 => x"2e9f38a9",
  1314 => x"ca048814",
  1315 => x"80f52d84",
  1316 => x"1508b4bc",
  1317 => x"53545285",
  1318 => x"f32d7184",
  1319 => x"29137008",
  1320 => x"5252a9ce",
  1321 => x"047351a8",
  1322 => x"992da9ca",
  1323 => x"04bd9008",
  1324 => x"8815082c",
  1325 => x"70810651",
  1326 => x"5271802e",
  1327 => x"8738b4c0",
  1328 => x"51a9c704",
  1329 => x"b4c45185",
  1330 => x"f32d8414",
  1331 => x"085185f3",
  1332 => x"2dbd9808",
  1333 => x"8105bd98",
  1334 => x"0c8c1454",
  1335 => x"a8d90402",
  1336 => x"90050d04",
  1337 => x"71bd940c",
  1338 => x"a8c92dbd",
  1339 => x"9808ff05",
  1340 => x"bd9c0c04",
  1341 => x"02ec050d",
  1342 => x"bd940855",
  1343 => x"80f851a7",
  1344 => x"b62db7e8",
  1345 => x"08812a70",
  1346 => x"81065152",
  1347 => x"719b3887",
  1348 => x"51a7b62d",
  1349 => x"b7e80881",
  1350 => x"2a708106",
  1351 => x"51527180",
  1352 => x"2eb138aa",
  1353 => x"a904a5ff",
  1354 => x"2d8751a7",
  1355 => x"b62db7e8",
  1356 => x"08f438aa",
  1357 => x"b904a5ff",
  1358 => x"2d80f851",
  1359 => x"a7b62db7",
  1360 => x"e808f338",
  1361 => x"b7e40881",
  1362 => x"3270b7e4",
  1363 => x"0c705252",
  1364 => x"84e52db7",
  1365 => x"e408a238",
  1366 => x"80da51a7",
  1367 => x"b62d81f5",
  1368 => x"51a7b62d",
  1369 => x"81f251a7",
  1370 => x"b62d81eb",
  1371 => x"51a7b62d",
  1372 => x"81f451a7",
  1373 => x"b62daebd",
  1374 => x"0481f551",
  1375 => x"a7b62db7",
  1376 => x"e808812a",
  1377 => x"70810651",
  1378 => x"5271802e",
  1379 => x"8f38bd9c",
  1380 => x"08527180",
  1381 => x"2e8638ff",
  1382 => x"12bd9c0c",
  1383 => x"81f251a7",
  1384 => x"b62db7e8",
  1385 => x"08812a70",
  1386 => x"81065152",
  1387 => x"71802e95",
  1388 => x"38bd9808",
  1389 => x"ff05bd9c",
  1390 => x"08545272",
  1391 => x"72258638",
  1392 => x"8113bd9c",
  1393 => x"0cbd9c08",
  1394 => x"70535473",
  1395 => x"802e8a38",
  1396 => x"8c15ff15",
  1397 => x"5555abcb",
  1398 => x"04820bb7",
  1399 => x"fc0c718f",
  1400 => x"06b7f80c",
  1401 => x"81eb51a7",
  1402 => x"b62db7e8",
  1403 => x"08812a70",
  1404 => x"81065152",
  1405 => x"71802ead",
  1406 => x"38740885",
  1407 => x"2e098106",
  1408 => x"a4388815",
  1409 => x"80f52dff",
  1410 => x"05527188",
  1411 => x"1681b72d",
  1412 => x"71982b52",
  1413 => x"71802588",
  1414 => x"38800b88",
  1415 => x"1681b72d",
  1416 => x"7451a899",
  1417 => x"2d81f451",
  1418 => x"a7b62db7",
  1419 => x"e808812a",
  1420 => x"70810651",
  1421 => x"5271802e",
  1422 => x"b3387408",
  1423 => x"852e0981",
  1424 => x"06aa3888",
  1425 => x"1580f52d",
  1426 => x"81055271",
  1427 => x"881681b7",
  1428 => x"2d7181ff",
  1429 => x"068b1680",
  1430 => x"f52d5452",
  1431 => x"72722787",
  1432 => x"38728816",
  1433 => x"81b72d74",
  1434 => x"51a8992d",
  1435 => x"80da51a7",
  1436 => x"b62db7e8",
  1437 => x"08812a70",
  1438 => x"81065152",
  1439 => x"71802e80",
  1440 => x"fb38bd94",
  1441 => x"08bd9c08",
  1442 => x"55537380",
  1443 => x"2e8a388c",
  1444 => x"13ff1555",
  1445 => x"53ad8a04",
  1446 => x"72085271",
  1447 => x"822ea638",
  1448 => x"71822689",
  1449 => x"3871812e",
  1450 => x"a538adfc",
  1451 => x"0471832e",
  1452 => x"ad387184",
  1453 => x"2e098106",
  1454 => x"80c23888",
  1455 => x"130851a9",
  1456 => x"e42dadfc",
  1457 => x"04881308",
  1458 => x"52712dad",
  1459 => x"fc04810b",
  1460 => x"8814082b",
  1461 => x"bd900832",
  1462 => x"bd900cad",
  1463 => x"f9048813",
  1464 => x"80f52d81",
  1465 => x"058b1480",
  1466 => x"f52d5354",
  1467 => x"71742483",
  1468 => x"38805473",
  1469 => x"881481b7",
  1470 => x"2da8c92d",
  1471 => x"8054800b",
  1472 => x"b7fc0c73",
  1473 => x"8f06b7f8",
  1474 => x"0ca05273",
  1475 => x"bd9c082e",
  1476 => x"09810698",
  1477 => x"38bd9808",
  1478 => x"ff057432",
  1479 => x"70098105",
  1480 => x"7072079f",
  1481 => x"2a917131",
  1482 => x"51515353",
  1483 => x"715182ee",
  1484 => x"2d811454",
  1485 => x"8e7425c6",
  1486 => x"38b7e408",
  1487 => x"5271b7e8",
  1488 => x"0c029405",
  1489 => x"0d040000",
  1490 => x"00ffffff",
  1491 => x"ff00ffff",
  1492 => x"ffff00ff",
  1493 => x"ffffff00",
  1494 => x"52657365",
  1495 => x"74000000",
  1496 => x"53617665",
  1497 => x"20616e64",
  1498 => x"20526573",
  1499 => x"65740000",
  1500 => x"4f707469",
  1501 => x"6f6e7320",
  1502 => x"10000000",
  1503 => x"536f756e",
  1504 => x"64201000",
  1505 => x"54757262",
  1506 => x"6f000000",
  1507 => x"4d6f7573",
  1508 => x"6520656d",
  1509 => x"756c6174",
  1510 => x"696f6e00",
  1511 => x"45786974",
  1512 => x"00000000",
  1513 => x"4d617374",
  1514 => x"65720000",
  1515 => x"4f504c4c",
  1516 => x"00000000",
  1517 => x"53434300",
  1518 => x"50534700",
  1519 => x"4261636b",
  1520 => x"00000000",
  1521 => x"5363616e",
  1522 => x"6c696e65",
  1523 => x"73000000",
  1524 => x"53442043",
  1525 => x"61726400",
  1526 => x"4a617061",
  1527 => x"6e657365",
  1528 => x"206b6579",
  1529 => x"206c6179",
  1530 => x"6f757400",
  1531 => x"32303438",
  1532 => x"4b422052",
  1533 => x"414d0000",
  1534 => x"34303936",
  1535 => x"4b422052",
  1536 => x"414d0000",
  1537 => x"536c323a",
  1538 => x"204e6f6e",
  1539 => x"65000000",
  1540 => x"536c323a",
  1541 => x"20455345",
  1542 => x"2d534343",
  1543 => x"20314d42",
  1544 => x"2f534343",
  1545 => x"2d490000",
  1546 => x"536c323a",
  1547 => x"20455345",
  1548 => x"2d52414d",
  1549 => x"20314d42",
  1550 => x"2f415343",
  1551 => x"49493800",
  1552 => x"536c323a",
  1553 => x"20455345",
  1554 => x"2d52414d",
  1555 => x"20314d42",
  1556 => x"2f415343",
  1557 => x"49493136",
  1558 => x"00000000",
  1559 => x"536c313a",
  1560 => x"204e6f6e",
  1561 => x"65000000",
  1562 => x"536c313a",
  1563 => x"20455345",
  1564 => x"2d534343",
  1565 => x"20314d42",
  1566 => x"2f534343",
  1567 => x"2d490000",
  1568 => x"536c313a",
  1569 => x"204d6567",
  1570 => x"6152414d",
  1571 => x"00000000",
  1572 => x"56474120",
  1573 => x"2d203331",
  1574 => x"4b487a2c",
  1575 => x"20363048",
  1576 => x"7a000000",
  1577 => x"56474120",
  1578 => x"2d203331",
  1579 => x"4b487a2c",
  1580 => x"20353048",
  1581 => x"7a000000",
  1582 => x"5456202d",
  1583 => x"20343830",
  1584 => x"692c2036",
  1585 => x"30487a00",
  1586 => x"496e6974",
  1587 => x"69616c69",
  1588 => x"7a696e67",
  1589 => x"20534420",
  1590 => x"63617264",
  1591 => x"0a000000",
  1592 => x"53444843",
  1593 => x"206e6f74",
  1594 => x"20737570",
  1595 => x"706f7274",
  1596 => x"65643b00",
  1597 => x"46617433",
  1598 => x"32206e6f",
  1599 => x"74207375",
  1600 => x"70706f72",
  1601 => x"7465643b",
  1602 => x"00000000",
  1603 => x"0a646973",
  1604 => x"61626c69",
  1605 => x"6e672053",
  1606 => x"44206361",
  1607 => x"72640a10",
  1608 => x"204f4b0a",
  1609 => x"00000000",
  1610 => x"4f434d53",
  1611 => x"58202020",
  1612 => x"43464700",
  1613 => x"54727969",
  1614 => x"6e67204d",
  1615 => x"53583342",
  1616 => x"494f532e",
  1617 => x"5359530a",
  1618 => x"00000000",
  1619 => x"4d535833",
  1620 => x"42494f53",
  1621 => x"53595300",
  1622 => x"54727969",
  1623 => x"6e672042",
  1624 => x"494f535f",
  1625 => x"4d32502e",
  1626 => x"524f4d0a",
  1627 => x"00000000",
  1628 => x"42494f53",
  1629 => x"5f4d3250",
  1630 => x"524f4d00",
  1631 => x"4c6f6164",
  1632 => x"696e6720",
  1633 => x"42494f53",
  1634 => x"0a000000",
  1635 => x"52656164",
  1636 => x"20666169",
  1637 => x"6c65640a",
  1638 => x"00000000",
  1639 => x"4c6f6164",
  1640 => x"696e6720",
  1641 => x"42494f53",
  1642 => x"20666169",
  1643 => x"6c65640a",
  1644 => x"00000000",
  1645 => x"4d425220",
  1646 => x"6661696c",
  1647 => x"0a000000",
  1648 => x"46415431",
  1649 => x"36202020",
  1650 => x"00000000",
  1651 => x"46415433",
  1652 => x"32202020",
  1653 => x"00000000",
  1654 => x"4e6f2070",
  1655 => x"61727469",
  1656 => x"74696f6e",
  1657 => x"20736967",
  1658 => x"0a000000",
  1659 => x"42616420",
  1660 => x"70617274",
  1661 => x"0a000000",
  1662 => x"53444843",
  1663 => x"20657272",
  1664 => x"6f72210a",
  1665 => x"00000000",
  1666 => x"53442069",
  1667 => x"6e69742e",
  1668 => x"2e2e0a00",
  1669 => x"53442063",
  1670 => x"61726420",
  1671 => x"72657365",
  1672 => x"74206661",
  1673 => x"696c6564",
  1674 => x"210a0000",
  1675 => x"57726974",
  1676 => x"65206661",
  1677 => x"696c6564",
  1678 => x"0a000000",
  1679 => x"16200000",
  1680 => x"14200000",
  1681 => x"15200000",
  1682 => x"00000002",
  1683 => x"00000002",
  1684 => x"00001758",
  1685 => x"0000067c",
  1686 => x"00000002",
  1687 => x"00001760",
  1688 => x"0000066e",
  1689 => x"00000004",
  1690 => x"00001770",
  1691 => x"00001af4",
  1692 => x"00000004",
  1693 => x"0000177c",
  1694 => x"00001aac",
  1695 => x"00000001",
  1696 => x"00001784",
  1697 => x"00000007",
  1698 => x"00000001",
  1699 => x"0000178c",
  1700 => x"0000000a",
  1701 => x"00000002",
  1702 => x"0000179c",
  1703 => x"00001406",
  1704 => x"00000000",
  1705 => x"00000000",
  1706 => x"00000000",
  1707 => x"00000005",
  1708 => x"000017a4",
  1709 => x"00000007",
  1710 => x"00000005",
  1711 => x"000017ac",
  1712 => x"00000007",
  1713 => x"00000005",
  1714 => x"000017b4",
  1715 => x"00000007",
  1716 => x"00000005",
  1717 => x"000017b8",
  1718 => x"00000007",
  1719 => x"00000004",
  1720 => x"000017bc",
  1721 => x"00001a4c",
  1722 => x"00000000",
  1723 => x"00000000",
  1724 => x"00000000",
  1725 => x"00000003",
  1726 => x"00001b84",
  1727 => x"00000003",
  1728 => x"00000001",
  1729 => x"000017c4",
  1730 => x"0000000b",
  1731 => x"00000001",
  1732 => x"000017d0",
  1733 => x"00000002",
  1734 => x"00000003",
  1735 => x"00001b78",
  1736 => x"00000003",
  1737 => x"00000003",
  1738 => x"00001b68",
  1739 => x"00000004",
  1740 => x"00000001",
  1741 => x"000017d8",
  1742 => x"00000006",
  1743 => x"00000003",
  1744 => x"00001b60",
  1745 => x"00000002",
  1746 => x"00000004",
  1747 => x"000017bc",
  1748 => x"00001a4c",
  1749 => x"00000000",
  1750 => x"00000000",
  1751 => x"00000000",
  1752 => x"000017ec",
  1753 => x"000017f8",
  1754 => x"00001804",
  1755 => x"00001810",
  1756 => x"00001828",
  1757 => x"00001840",
  1758 => x"0000185c",
  1759 => x"00001868",
  1760 => x"00001880",
  1761 => x"00001890",
  1762 => x"000018a4",
  1763 => x"000018b8",
  1764 => x"00000003",
  1765 => x"00000000",
  1766 => x"00000000",
  1767 => x"00000000",
  1768 => x"00000000",
  1769 => x"00000000",
  1770 => x"00000000",
  1771 => x"00000000",
  1772 => x"00000000",
  1773 => x"00000000",
  1774 => x"00000000",
  1775 => x"00000000",
  1776 => x"00000000",
  1777 => x"00000000",
  1778 => x"00000000",
  1779 => x"00000000",
  1780 => x"00000000",
  1781 => x"00000000",
  1782 => x"00000000",
  1783 => x"00000000",
  1784 => x"00000000",
  1785 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

