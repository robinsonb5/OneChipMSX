-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b0bb7",
     9 => x"c8080b0b",
    10 => x"0bb7cc08",
    11 => x"0b0b0bb7",
    12 => x"d0080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"b7d00c0b",
    16 => x"0b0bb7cc",
    17 => x"0c0b0b0b",
    18 => x"b7c80c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0baea4",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"b7c870bd",
    57 => x"80278b38",
    58 => x"80717084",
    59 => x"05530c81",
    60 => x"e2048c51",
    61 => x"8d8d0402",
    62 => x"fc050df8",
    63 => x"80518f0b",
    64 => x"b7d80c9f",
    65 => x"0bb7dc0c",
    66 => x"a0717081",
    67 => x"055334b7",
    68 => x"dc08ff05",
    69 => x"b7dc0cb7",
    70 => x"dc088025",
    71 => x"eb38b7d8",
    72 => x"08ff05b7",
    73 => x"d80cb7d8",
    74 => x"088025d7",
    75 => x"38028405",
    76 => x"0d0402f0",
    77 => x"050df880",
    78 => x"53f8a054",
    79 => x"83bf5273",
    80 => x"70810555",
    81 => x"33517073",
    82 => x"70810555",
    83 => x"34ff1252",
    84 => x"718025eb",
    85 => x"38fbc053",
    86 => x"9f52a073",
    87 => x"70810555",
    88 => x"34ff1252",
    89 => x"718025f2",
    90 => x"38029005",
    91 => x"0d0402f4",
    92 => x"050d7453",
    93 => x"8e0bb7d8",
    94 => x"08258f38",
    95 => x"82b22db7",
    96 => x"d808ff05",
    97 => x"b7d80c82",
    98 => x"f404b7d8",
    99 => x"08b7dc08",
   100 => x"5351728a",
   101 => x"2e098106",
   102 => x"b7387151",
   103 => x"719f24a0",
   104 => x"38b7d808",
   105 => x"a02911f8",
   106 => x"80115151",
   107 => x"a07134b7",
   108 => x"dc088105",
   109 => x"b7dc0cb7",
   110 => x"dc08519f",
   111 => x"7125e238",
   112 => x"800bb7dc",
   113 => x"0cb7d808",
   114 => x"8105b7d8",
   115 => x"0c83e404",
   116 => x"70a02912",
   117 => x"f8801151",
   118 => x"51727134",
   119 => x"b7dc0881",
   120 => x"05b7dc0c",
   121 => x"b7dc08a0",
   122 => x"2e098106",
   123 => x"8e38800b",
   124 => x"b7dc0cb7",
   125 => x"d8088105",
   126 => x"b7d80c02",
   127 => x"8c050d04",
   128 => x"02e8050d",
   129 => x"77795656",
   130 => x"880bfc16",
   131 => x"77712c8f",
   132 => x"06545254",
   133 => x"80537272",
   134 => x"25953871",
   135 => x"53fbe014",
   136 => x"51877134",
   137 => x"8114ff14",
   138 => x"545472f1",
   139 => x"387153f9",
   140 => x"1576712c",
   141 => x"87065351",
   142 => x"71802e8b",
   143 => x"38fbe014",
   144 => x"51717134",
   145 => x"81145472",
   146 => x"8e249538",
   147 => x"8f733153",
   148 => x"fbe01451",
   149 => x"a0713481",
   150 => x"14ff1454",
   151 => x"5472f138",
   152 => x"0298050d",
   153 => x"0402ec05",
   154 => x"0d800bb7",
   155 => x"e00cf68c",
   156 => x"08f69008",
   157 => x"71882c56",
   158 => x"5481ff06",
   159 => x"52737225",
   160 => x"88387154",
   161 => x"820bb7e0",
   162 => x"0c72882c",
   163 => x"7381ff06",
   164 => x"54557473",
   165 => x"258b3872",
   166 => x"b7e00884",
   167 => x"07b7e00c",
   168 => x"5573842b",
   169 => x"86a07125",
   170 => x"83713170",
   171 => x"0b0b0bb4",
   172 => x"a40c8171",
   173 => x"2bff05f6",
   174 => x"880cfecc",
   175 => x"13ff122c",
   176 => x"788829ff",
   177 => x"94057081",
   178 => x"2cb7e008",
   179 => x"52585255",
   180 => x"51525476",
   181 => x"802e8538",
   182 => x"70810751",
   183 => x"70f6940c",
   184 => x"71098105",
   185 => x"f6800c72",
   186 => x"098105f6",
   187 => x"840c0294",
   188 => x"050d0402",
   189 => x"f4050d74",
   190 => x"53727081",
   191 => x"055480f5",
   192 => x"2d527180",
   193 => x"2e893871",
   194 => x"5182ee2d",
   195 => x"85f90402",
   196 => x"8c050d04",
   197 => x"02f8050d",
   198 => x"a5da2d80",
   199 => x"da51a791",
   200 => x"2db7c808",
   201 => x"812a7081",
   202 => x"06515271",
   203 => x"802ee938",
   204 => x"0288050d",
   205 => x"0402f405",
   206 => x"0dbcf008",
   207 => x"99c406b6",
   208 => x"a00b80f5",
   209 => x"2d525270",
   210 => x"802e8638",
   211 => x"71848007",
   212 => x"52b5d80b",
   213 => x"80f52d72",
   214 => x"07b5fc0b",
   215 => x"80f52d70",
   216 => x"812a7081",
   217 => x"06515354",
   218 => x"5270802e",
   219 => x"86387182",
   220 => x"80075272",
   221 => x"81065170",
   222 => x"802e8538",
   223 => x"71880752",
   224 => x"b6880b80",
   225 => x"f52d7084",
   226 => x"2b730781",
   227 => x"8432b7c8",
   228 => x"0c51028c",
   229 => x"050d0402",
   230 => x"f4050d74",
   231 => x"70818432",
   232 => x"bcf00c70",
   233 => x"83065253",
   234 => x"70b5d00b",
   235 => x"880581b7",
   236 => x"2d72892a",
   237 => x"70810651",
   238 => x"5170b6a0",
   239 => x"0b81b72d",
   240 => x"72832a81",
   241 => x"0673882a",
   242 => x"70810651",
   243 => x"52527080",
   244 => x"2e853871",
   245 => x"82075271",
   246 => x"b5fc0b81",
   247 => x"b72d7284",
   248 => x"2c708306",
   249 => x"515170b6",
   250 => x"880b81b7",
   251 => x"2d70b7c8",
   252 => x"0c028c05",
   253 => x"0d0402f4",
   254 => x"050db588",
   255 => x"0b881180",
   256 => x"f52d8c12",
   257 => x"881180f5",
   258 => x"2d70842b",
   259 => x"73078c13",
   260 => x"881180f5",
   261 => x"2d70882b",
   262 => x"73079413",
   263 => x"80f52d70",
   264 => x"8c2b7207",
   265 => x"b7c80c53",
   266 => x"53535353",
   267 => x"56525351",
   268 => x"028c050d",
   269 => x"0402f405",
   270 => x"0d74b588",
   271 => x"71870655",
   272 => x"53517288",
   273 => x"1381b72d",
   274 => x"8c127184",
   275 => x"2c708706",
   276 => x"55525272",
   277 => x"881381b7",
   278 => x"2d8c1271",
   279 => x"842c7087",
   280 => x"06555252",
   281 => x"72881381",
   282 => x"b72d7084",
   283 => x"2c708706",
   284 => x"51517094",
   285 => x"1381b72d",
   286 => x"028c050d",
   287 => x"0402d405",
   288 => x"0db1a451",
   289 => x"85f32d9d",
   290 => x"be2db7c8",
   291 => x"08802e83",
   292 => x"a23886b5",
   293 => x"2db7c808",
   294 => x"5390872d",
   295 => x"b7c80854",
   296 => x"b7c80880",
   297 => x"2e838e38",
   298 => x"a1c12db7",
   299 => x"c808802e",
   300 => x"8738b1bc",
   301 => x"5189c504",
   302 => x"99aa2db7",
   303 => x"c808802e",
   304 => x"a238b1d0",
   305 => x"5185f32d",
   306 => x"b1e85185",
   307 => x"f32d8694",
   308 => x"2d728407",
   309 => x"53810bfe",
   310 => x"c40c72fe",
   311 => x"c00c7251",
   312 => x"87972d84",
   313 => x"0bfec40c",
   314 => x"b28452b7",
   315 => x"e8519699",
   316 => x"2db7c808",
   317 => x"802e80e1",
   318 => x"387c802e",
   319 => x"af3872b7",
   320 => x"f40c87f6",
   321 => x"2db7c808",
   322 => x"b7f80cb7",
   323 => x"fc5480fd",
   324 => x"53807470",
   325 => x"8405560c",
   326 => x"ff135372",
   327 => x"8025f238",
   328 => x"b7f452b7",
   329 => x"e8519984",
   330 => x"2d8ad904",
   331 => x"b28452b7",
   332 => x"e8519699",
   333 => x"2db7c808",
   334 => x"802e9e38",
   335 => x"b7f452b7",
   336 => x"e85198de",
   337 => x"2db7f408",
   338 => x"b7f80852",
   339 => x"5388b52d",
   340 => x"72fec00c",
   341 => x"72518797",
   342 => x"2db29051",
   343 => x"85f32db2",
   344 => x"a852b7e8",
   345 => x"5196992d",
   346 => x"b7c80898",
   347 => x"38b2b451",
   348 => x"85f32db2",
   349 => x"cc52b7e8",
   350 => x"5196992d",
   351 => x"b7c80880",
   352 => x"2e81b038",
   353 => x"b2d85185",
   354 => x"f32db7ec",
   355 => x"08578077",
   356 => x"595a767a",
   357 => x"2e8b3881",
   358 => x"1a78812a",
   359 => x"595a77f7",
   360 => x"38f71a5a",
   361 => x"80772581",
   362 => x"80387952",
   363 => x"77518480",
   364 => x"2db7f452",
   365 => x"b7e85198",
   366 => x"de2db7c8",
   367 => x"0853b7c8",
   368 => x"08802e80",
   369 => x"c938b7f4",
   370 => x"5b80598b",
   371 => x"fb047a70",
   372 => x"84055c08",
   373 => x"7081ff06",
   374 => x"71882c70",
   375 => x"81ff0673",
   376 => x"902c7081",
   377 => x"ff067598",
   378 => x"2afec80c",
   379 => x"fec80c58",
   380 => x"fec80c57",
   381 => x"fec80c84",
   382 => x"1a5a5376",
   383 => x"53848077",
   384 => x"25843884",
   385 => x"80537279",
   386 => x"24c4388c",
   387 => x"9904b2e8",
   388 => x"5185f32d",
   389 => x"72548cb5",
   390 => x"04b7e851",
   391 => x"98b12dfc",
   392 => x"80178119",
   393 => x"59578ba4",
   394 => x"04820bfe",
   395 => x"c40c8154",
   396 => x"8cb50480",
   397 => x"5473b7c8",
   398 => x"0c02ac05",
   399 => x"0d0402f8",
   400 => x"050da7e1",
   401 => x"2d81f72d",
   402 => x"815184e5",
   403 => x"2dfec452",
   404 => x"81720ca5",
   405 => x"a12da5a1",
   406 => x"2d84720c",
   407 => x"735188fd",
   408 => x"2db4a851",
   409 => x"a9bf2d80",
   410 => x"5184e52d",
   411 => x"0288050d",
   412 => x"0402fc05",
   413 => x"0d81518c",
   414 => x"be2d0284",
   415 => x"050d0402",
   416 => x"fc050d80",
   417 => x"518cbe2d",
   418 => x"0284050d",
   419 => x"0402ec05",
   420 => x"0d84b851",
   421 => x"87972d81",
   422 => x"0bfec40c",
   423 => x"84b80bfe",
   424 => x"c00c840b",
   425 => x"fec40c83",
   426 => x"0bfecc0c",
   427 => x"a5bc2da7",
   428 => x"d52da5a1",
   429 => x"2da5a12d",
   430 => x"81f72d81",
   431 => x"5184e52d",
   432 => x"a5a12da5",
   433 => x"a12d8151",
   434 => x"84e52d80",
   435 => x"5188fd2d",
   436 => x"b7c80880",
   437 => x"2e81dd38",
   438 => x"805184e5",
   439 => x"2db4a851",
   440 => x"a9bf2dbc",
   441 => x"d8080970",
   442 => x"8306fecc",
   443 => x"0c52bcd0",
   444 => x"088938bc",
   445 => x"d408802e",
   446 => x"80e238fe",
   447 => x"d0087081",
   448 => x"06515271",
   449 => x"802e80d4",
   450 => x"38a7db2d",
   451 => x"bcd00870",
   452 => x"bcd40870",
   453 => x"57555652",
   454 => x"80ff7225",
   455 => x"843880ff",
   456 => x"5280ff73",
   457 => x"25843880",
   458 => x"ff5371ff",
   459 => x"80258438",
   460 => x"ff805272",
   461 => x"ff802584",
   462 => x"38ff8053",
   463 => x"747231bc",
   464 => x"d00c7373",
   465 => x"31bcd40c",
   466 => x"a7d52d71",
   467 => x"882b83fe",
   468 => x"80067381",
   469 => x"ff067107",
   470 => x"fed00c52",
   471 => x"a5da2da9",
   472 => x"cf2db7c8",
   473 => x"085386b5",
   474 => x"2db7c808",
   475 => x"fec00c87",
   476 => x"f62db7c8",
   477 => x"08fed40c",
   478 => x"86b52db7",
   479 => x"c808b7e4",
   480 => x"082e9c38",
   481 => x"b7c808b7",
   482 => x"e40c8452",
   483 => x"725184e5",
   484 => x"2da5a12d",
   485 => x"a5a12dff",
   486 => x"12527180",
   487 => x"25ee3872",
   488 => x"802e8938",
   489 => x"8a0bfec4",
   490 => x"0c8de304",
   491 => x"820bfec4",
   492 => x"0c8de304",
   493 => x"b2f85185",
   494 => x"f32d820b",
   495 => x"fec40c80",
   496 => x"0bb7c80c",
   497 => x"0294050d",
   498 => x"0402e805",
   499 => x"0d77797b",
   500 => x"58555580",
   501 => x"53727625",
   502 => x"a3387470",
   503 => x"81055680",
   504 => x"f52d7470",
   505 => x"81055680",
   506 => x"f52d5252",
   507 => x"71712e86",
   508 => x"3881518f",
   509 => x"fe048113",
   510 => x"538fd504",
   511 => x"805170b7",
   512 => x"c80c0298",
   513 => x"050d0402",
   514 => x"d8050d80",
   515 => x"0bbbfc0c",
   516 => x"b7f45280",
   517 => x"51a0a62d",
   518 => x"b7c80854",
   519 => x"b7c8088c",
   520 => x"38b39051",
   521 => x"85f32d73",
   522 => x"5595a204",
   523 => x"8056810b",
   524 => x"bca00c88",
   525 => x"53b39c52",
   526 => x"b8aa518f",
   527 => x"c92db7c8",
   528 => x"08762e09",
   529 => x"81068738",
   530 => x"b7c808bc",
   531 => x"a00c8853",
   532 => x"b3a852b8",
   533 => x"c6518fc9",
   534 => x"2db7c808",
   535 => x"8738b7c8",
   536 => x"08bca00c",
   537 => x"bca00880",
   538 => x"2e80f638",
   539 => x"bbba0b80",
   540 => x"f52dbbbb",
   541 => x"0b80f52d",
   542 => x"71982b71",
   543 => x"902b07bb",
   544 => x"bc0b80f5",
   545 => x"2d70882b",
   546 => x"7207bbbd",
   547 => x"0b80f52d",
   548 => x"7107bbf2",
   549 => x"0b80f52d",
   550 => x"bbf30b80",
   551 => x"f52d7188",
   552 => x"2b07535f",
   553 => x"54525a56",
   554 => x"57557381",
   555 => x"abaa2e09",
   556 => x"81068d38",
   557 => x"7551a1c8",
   558 => x"2db7c808",
   559 => x"5691cd04",
   560 => x"7382d4d5",
   561 => x"2e8738b3",
   562 => x"b451928e",
   563 => x"04b7f452",
   564 => x"7551a0a6",
   565 => x"2db7c808",
   566 => x"55b7c808",
   567 => x"802e83c2",
   568 => x"388853b3",
   569 => x"a852b8c6",
   570 => x"518fc92d",
   571 => x"b7c80889",
   572 => x"38810bbb",
   573 => x"fc0c9294",
   574 => x"048853b3",
   575 => x"9c52b8aa",
   576 => x"518fc92d",
   577 => x"b7c80880",
   578 => x"2e8a38b3",
   579 => x"c85185f3",
   580 => x"2d92ee04",
   581 => x"bbf20b80",
   582 => x"f52d5473",
   583 => x"80d52e09",
   584 => x"810680ca",
   585 => x"38bbf30b",
   586 => x"80f52d54",
   587 => x"7381aa2e",
   588 => x"098106ba",
   589 => x"38800bb7",
   590 => x"f40b80f5",
   591 => x"2d565474",
   592 => x"81e92e83",
   593 => x"38815474",
   594 => x"81eb2e8c",
   595 => x"38805573",
   596 => x"752e0981",
   597 => x"0682cb38",
   598 => x"b7ff0b80",
   599 => x"f52d5574",
   600 => x"8d38b880",
   601 => x"0b80f52d",
   602 => x"5473822e",
   603 => x"86388055",
   604 => x"95a204b8",
   605 => x"810b80f5",
   606 => x"2d70bbf4",
   607 => x"0cff05bb",
   608 => x"f80cb882",
   609 => x"0b80f52d",
   610 => x"b8830b80",
   611 => x"f52d5876",
   612 => x"05778280",
   613 => x"290570bc",
   614 => x"800cb884",
   615 => x"0b80f52d",
   616 => x"70bc940c",
   617 => x"bbfc0859",
   618 => x"57587680",
   619 => x"2e81a338",
   620 => x"8853b3a8",
   621 => x"52b8c651",
   622 => x"8fc92db7",
   623 => x"c80881e2",
   624 => x"38bbf408",
   625 => x"70842bbc",
   626 => x"980c70bc",
   627 => x"900cb899",
   628 => x"0b80f52d",
   629 => x"b8980b80",
   630 => x"f52d7182",
   631 => x"802905b8",
   632 => x"9a0b80f5",
   633 => x"2d708480",
   634 => x"802912b8",
   635 => x"9b0b80f5",
   636 => x"2d708180",
   637 => x"0a291270",
   638 => x"bc9c0cbc",
   639 => x"94087129",
   640 => x"bc800805",
   641 => x"70bc840c",
   642 => x"b8a10b80",
   643 => x"f52db8a0",
   644 => x"0b80f52d",
   645 => x"71828029",
   646 => x"05b8a20b",
   647 => x"80f52d70",
   648 => x"84808029",
   649 => x"12b8a30b",
   650 => x"80f52d70",
   651 => x"982b81f0",
   652 => x"0a067205",
   653 => x"70bc880c",
   654 => x"fe117e29",
   655 => x"7705bc8c",
   656 => x"0c525952",
   657 => x"43545e51",
   658 => x"5259525d",
   659 => x"57595795",
   660 => x"a004b886",
   661 => x"0b80f52d",
   662 => x"b8850b80",
   663 => x"f52d7182",
   664 => x"80290570",
   665 => x"bc980c70",
   666 => x"a02983ff",
   667 => x"0570892a",
   668 => x"70bc900c",
   669 => x"b88b0b80",
   670 => x"f52db88a",
   671 => x"0b80f52d",
   672 => x"71828029",
   673 => x"0570bc9c",
   674 => x"0c7b7129",
   675 => x"1e70bc8c",
   676 => x"0c7dbc88",
   677 => x"0c7305bc",
   678 => x"840c555e",
   679 => x"51515555",
   680 => x"815574b7",
   681 => x"c80c02a8",
   682 => x"050d0402",
   683 => x"ec050d76",
   684 => x"70872c71",
   685 => x"80ff0655",
   686 => x"5654bbfc",
   687 => x"088a3873",
   688 => x"882c7481",
   689 => x"ff065455",
   690 => x"b7f452bc",
   691 => x"80081551",
   692 => x"a0a62db7",
   693 => x"c80854b7",
   694 => x"c808802e",
   695 => x"b338bbfc",
   696 => x"08802e98",
   697 => x"38728429",
   698 => x"b7f40570",
   699 => x"085253a1",
   700 => x"c82db7c8",
   701 => x"08f00a06",
   702 => x"53968e04",
   703 => x"7210b7f4",
   704 => x"057080e0",
   705 => x"2d5253a1",
   706 => x"f82db7c8",
   707 => x"08537254",
   708 => x"73b7c80c",
   709 => x"0294050d",
   710 => x"0402c805",
   711 => x"0d7f615f",
   712 => x"5b800bbc",
   713 => x"8808bc8c",
   714 => x"08595d56",
   715 => x"bbfc0876",
   716 => x"2e8a38bb",
   717 => x"f408842b",
   718 => x"5896c204",
   719 => x"bc900884",
   720 => x"2b588059",
   721 => x"78782781",
   722 => x"a938788f",
   723 => x"06a01757",
   724 => x"54738f38",
   725 => x"b7f45276",
   726 => x"51811757",
   727 => x"a0a62db7",
   728 => x"f4568076",
   729 => x"80f52d56",
   730 => x"5474742e",
   731 => x"83388154",
   732 => x"7481e52e",
   733 => x"80f63881",
   734 => x"70750655",
   735 => x"5d73802e",
   736 => x"80ea388b",
   737 => x"1680f52d",
   738 => x"98065a79",
   739 => x"80de388b",
   740 => x"537d5275",
   741 => x"518fc92d",
   742 => x"b7c80880",
   743 => x"cf389c16",
   744 => x"0851a1c8",
   745 => x"2db7c808",
   746 => x"841c0c9a",
   747 => x"1680e02d",
   748 => x"51a1f82d",
   749 => x"b7c808b7",
   750 => x"c808881d",
   751 => x"0cb7c808",
   752 => x"5555bbfc",
   753 => x"08802e98",
   754 => x"38941680",
   755 => x"e02d51a1",
   756 => x"f82db7c8",
   757 => x"08902b83",
   758 => x"fff00a06",
   759 => x"70165154",
   760 => x"73881c0c",
   761 => x"797b0c7c",
   762 => x"5498a804",
   763 => x"81195996",
   764 => x"c404bbfc",
   765 => x"08802eae",
   766 => x"387b5195",
   767 => x"ab2db7c8",
   768 => x"08b7c808",
   769 => x"80ffffff",
   770 => x"f806555c",
   771 => x"7380ffff",
   772 => x"fff82e92",
   773 => x"38b7c808",
   774 => x"fe05bbf4",
   775 => x"0829bc84",
   776 => x"08055796",
   777 => x"c2048054",
   778 => x"73b7c80c",
   779 => x"02b8050d",
   780 => x"0402f405",
   781 => x"0d747008",
   782 => x"8105710c",
   783 => x"7008bbf8",
   784 => x"08065353",
   785 => x"718e3888",
   786 => x"13085195",
   787 => x"ab2db7c8",
   788 => x"0888140c",
   789 => x"810bb7c8",
   790 => x"0c028c05",
   791 => x"0d0402f0",
   792 => x"050d7588",
   793 => x"1108fe05",
   794 => x"bbf40829",
   795 => x"bc840811",
   796 => x"7208bbf8",
   797 => x"08060579",
   798 => x"55535454",
   799 => x"a0a62d02",
   800 => x"90050d04",
   801 => x"02f0050d",
   802 => x"75881108",
   803 => x"fe05bbf4",
   804 => x"0829bc84",
   805 => x"08117208",
   806 => x"bbf80806",
   807 => x"05795553",
   808 => x"54549ee6",
   809 => x"2d029005",
   810 => x"0d04bbfc",
   811 => x"08b7c80c",
   812 => x"0402f405",
   813 => x"0dd45281",
   814 => x"ff720c71",
   815 => x"085381ff",
   816 => x"720c7288",
   817 => x"2b83fe80",
   818 => x"06720870",
   819 => x"81ff0651",
   820 => x"525381ff",
   821 => x"720c7271",
   822 => x"07882b72",
   823 => x"087081ff",
   824 => x"06515253",
   825 => x"81ff720c",
   826 => x"72710788",
   827 => x"2b720870",
   828 => x"81ff0672",
   829 => x"07b7c80c",
   830 => x"5253028c",
   831 => x"050d0402",
   832 => x"f4050d74",
   833 => x"767181ff",
   834 => x"06d40c53",
   835 => x"53bca408",
   836 => x"85387189",
   837 => x"2b527198",
   838 => x"2ad40c71",
   839 => x"902a7081",
   840 => x"ff06d40c",
   841 => x"5171882a",
   842 => x"7081ff06",
   843 => x"d40c5171",
   844 => x"81ff06d4",
   845 => x"0c72902a",
   846 => x"7081ff06",
   847 => x"d40c51d4",
   848 => x"087081ff",
   849 => x"06515182",
   850 => x"b8bf5270",
   851 => x"81ff2e09",
   852 => x"81069438",
   853 => x"81ff0bd4",
   854 => x"0cd40870",
   855 => x"81ff06ff",
   856 => x"14545151",
   857 => x"71e53870",
   858 => x"b7c80c02",
   859 => x"8c050d04",
   860 => x"02fc050d",
   861 => x"81c75181",
   862 => x"ff0bd40c",
   863 => x"ff115170",
   864 => x"8025f438",
   865 => x"0284050d",
   866 => x"0402f005",
   867 => x"0d9af02d",
   868 => x"8fcf5380",
   869 => x"5287fc80",
   870 => x"f75199ff",
   871 => x"2db7c808",
   872 => x"54b7c808",
   873 => x"812e0981",
   874 => x"06a33881",
   875 => x"ff0bd40c",
   876 => x"820a5284",
   877 => x"9c80e951",
   878 => x"99ff2db7",
   879 => x"c8088b38",
   880 => x"81ff0bd4",
   881 => x"0c73539b",
   882 => x"d3049af0",
   883 => x"2dff1353",
   884 => x"72c13872",
   885 => x"b7c80c02",
   886 => x"90050d04",
   887 => x"02f4050d",
   888 => x"81ff0bd4",
   889 => x"0c935380",
   890 => x"5287fc80",
   891 => x"c15199ff",
   892 => x"2db7c808",
   893 => x"8b3881ff",
   894 => x"0bd40c81",
   895 => x"539c8904",
   896 => x"9af02dff",
   897 => x"135372df",
   898 => x"3872b7c8",
   899 => x"0c028c05",
   900 => x"0d0402f0",
   901 => x"050d9af0",
   902 => x"2d83aa52",
   903 => x"849c80c8",
   904 => x"5199ff2d",
   905 => x"b7c80881",
   906 => x"2e098106",
   907 => x"923899b1",
   908 => x"2db7c808",
   909 => x"83ffff06",
   910 => x"537283aa",
   911 => x"2e97389b",
   912 => x"dc2d9cd0",
   913 => x"0481549d",
   914 => x"b504b3d4",
   915 => x"5185f32d",
   916 => x"80549db5",
   917 => x"0481ff0b",
   918 => x"d40cb153",
   919 => x"9b892db7",
   920 => x"c808802e",
   921 => x"80c03880",
   922 => x"5287fc80",
   923 => x"fa5199ff",
   924 => x"2db7c808",
   925 => x"b13881ff",
   926 => x"0bd40cd4",
   927 => x"085381ff",
   928 => x"0bd40c81",
   929 => x"ff0bd40c",
   930 => x"81ff0bd4",
   931 => x"0c81ff0b",
   932 => x"d40c7286",
   933 => x"2a708106",
   934 => x"b7c80856",
   935 => x"51537280",
   936 => x"2e93389c",
   937 => x"c5047282",
   938 => x"2eff9f38",
   939 => x"ff135372",
   940 => x"ffaa3872",
   941 => x"5473b7c8",
   942 => x"0c029005",
   943 => x"0d0402f0",
   944 => x"050d810b",
   945 => x"bca40c84",
   946 => x"54d00870",
   947 => x"8f2a7081",
   948 => x"06515153",
   949 => x"72f33872",
   950 => x"d00c9af0",
   951 => x"2db3e451",
   952 => x"85f32dd0",
   953 => x"08708f2a",
   954 => x"70810651",
   955 => x"515372f3",
   956 => x"38810bd0",
   957 => x"0cb15380",
   958 => x"5284d480",
   959 => x"c05199ff",
   960 => x"2db7c808",
   961 => x"812ea138",
   962 => x"72822e09",
   963 => x"81068c38",
   964 => x"b3f05185",
   965 => x"f32d8053",
   966 => x"9edd04ff",
   967 => x"135372d7",
   968 => x"38ff1454",
   969 => x"73ffa238",
   970 => x"9c922db7",
   971 => x"c808bca4",
   972 => x"0cb7c808",
   973 => x"8b388152",
   974 => x"87fc80d0",
   975 => x"5199ff2d",
   976 => x"81ff0bd4",
   977 => x"0cd00870",
   978 => x"8f2a7081",
   979 => x"06515153",
   980 => x"72f33872",
   981 => x"d00c81ff",
   982 => x"0bd40c81",
   983 => x"5372b7c8",
   984 => x"0c029005",
   985 => x"0d0402e8",
   986 => x"050d7856",
   987 => x"81ff0bd4",
   988 => x"0cd00870",
   989 => x"8f2a7081",
   990 => x"06515153",
   991 => x"72f33882",
   992 => x"810bd00c",
   993 => x"81ff0bd4",
   994 => x"0c775287",
   995 => x"fc80d851",
   996 => x"99ff2db7",
   997 => x"c808802e",
   998 => x"8c38b488",
   999 => x"5185f32d",
  1000 => x"8153a09d",
  1001 => x"0481ff0b",
  1002 => x"d40c81fe",
  1003 => x"0bd40c80",
  1004 => x"ff557570",
  1005 => x"84055708",
  1006 => x"70982ad4",
  1007 => x"0c70902c",
  1008 => x"7081ff06",
  1009 => x"d40c5470",
  1010 => x"882c7081",
  1011 => x"ff06d40c",
  1012 => x"547081ff",
  1013 => x"06d40c54",
  1014 => x"ff155574",
  1015 => x"8025d338",
  1016 => x"81ff0bd4",
  1017 => x"0c81ff0b",
  1018 => x"d40c81ff",
  1019 => x"0bd40c86",
  1020 => x"8da05481",
  1021 => x"ff0bd40c",
  1022 => x"d40881ff",
  1023 => x"06557487",
  1024 => x"38ff1454",
  1025 => x"73ed3881",
  1026 => x"ff0bd40c",
  1027 => x"d008708f",
  1028 => x"2a708106",
  1029 => x"51515372",
  1030 => x"f33872d0",
  1031 => x"0c72b7c8",
  1032 => x"0c029805",
  1033 => x"0d0402e8",
  1034 => x"050d7855",
  1035 => x"805681ff",
  1036 => x"0bd40cd0",
  1037 => x"08708f2a",
  1038 => x"70810651",
  1039 => x"515372f3",
  1040 => x"3882810b",
  1041 => x"d00c81ff",
  1042 => x"0bd40c77",
  1043 => x"5287fc80",
  1044 => x"d15199ff",
  1045 => x"2d80dbc6",
  1046 => x"df54b7c8",
  1047 => x"08802e8a",
  1048 => x"38b2e851",
  1049 => x"85f32da1",
  1050 => x"b80481ff",
  1051 => x"0bd40cd4",
  1052 => x"087081ff",
  1053 => x"06515372",
  1054 => x"81fe2e09",
  1055 => x"81069d38",
  1056 => x"80ff5399",
  1057 => x"b12db7c8",
  1058 => x"08757084",
  1059 => x"05570cff",
  1060 => x"13537280",
  1061 => x"25ed3881",
  1062 => x"56a1a204",
  1063 => x"ff145473",
  1064 => x"c93881ff",
  1065 => x"0bd40cd0",
  1066 => x"08708f2a",
  1067 => x"70810651",
  1068 => x"515372f3",
  1069 => x"3872d00c",
  1070 => x"75b7c80c",
  1071 => x"0298050d",
  1072 => x"04bca408",
  1073 => x"b7c80c04",
  1074 => x"02f4050d",
  1075 => x"7470882a",
  1076 => x"83fe8006",
  1077 => x"7072982a",
  1078 => x"0772882b",
  1079 => x"87fc8080",
  1080 => x"0673982b",
  1081 => x"81f00a06",
  1082 => x"71730707",
  1083 => x"b7c80c56",
  1084 => x"51535102",
  1085 => x"8c050d04",
  1086 => x"02f8050d",
  1087 => x"028e0580",
  1088 => x"f52d7488",
  1089 => x"2b077083",
  1090 => x"ffff06b7",
  1091 => x"c80c5102",
  1092 => x"88050d04",
  1093 => x"02fc050d",
  1094 => x"72518071",
  1095 => x"0c800b84",
  1096 => x"120c0284",
  1097 => x"050d0402",
  1098 => x"f0050d75",
  1099 => x"70088412",
  1100 => x"08535353",
  1101 => x"ff547171",
  1102 => x"2ea838a7",
  1103 => x"db2d8413",
  1104 => x"08708429",
  1105 => x"14881170",
  1106 => x"087081ff",
  1107 => x"06841808",
  1108 => x"81118706",
  1109 => x"841a0c53",
  1110 => x"51555151",
  1111 => x"51a7d52d",
  1112 => x"715473b7",
  1113 => x"c80c0290",
  1114 => x"050d0402",
  1115 => x"f0050da7",
  1116 => x"db2de008",
  1117 => x"e408718b",
  1118 => x"2a708106",
  1119 => x"51535552",
  1120 => x"70802e9d",
  1121 => x"38bca808",
  1122 => x"708429bc",
  1123 => x"b0057381",
  1124 => x"ff06710c",
  1125 => x"5151bca8",
  1126 => x"08811187",
  1127 => x"06bca80c",
  1128 => x"51738b2a",
  1129 => x"70810651",
  1130 => x"5170802e",
  1131 => x"818938b6",
  1132 => x"f8088429",
  1133 => x"bce00574",
  1134 => x"81ff0671",
  1135 => x"0c51b6f8",
  1136 => x"088105b6",
  1137 => x"f80c850b",
  1138 => x"b6f40cb6",
  1139 => x"f808b6f0",
  1140 => x"082e0981",
  1141 => x"06818638",
  1142 => x"800bb6f8",
  1143 => x"0cbce008",
  1144 => x"708306bc",
  1145 => x"d80c7085",
  1146 => x"2a708106",
  1147 => x"bcd40856",
  1148 => x"51525270",
  1149 => x"802e8e38",
  1150 => x"bce808fe",
  1151 => x"803213bc",
  1152 => x"d40ca48c",
  1153 => x"04bce808",
  1154 => x"13bcd40c",
  1155 => x"71842a70",
  1156 => x"8106bcd0",
  1157 => x"08545151",
  1158 => x"70802e90",
  1159 => x"38bce408",
  1160 => x"81ff3212",
  1161 => x"8105bcd0",
  1162 => x"0ca4dd04",
  1163 => x"71bce408",
  1164 => x"31bcd00c",
  1165 => x"a4dd04b6",
  1166 => x"f408ff05",
  1167 => x"b6f40cb6",
  1168 => x"f408ff2e",
  1169 => x"09810695",
  1170 => x"38b6f808",
  1171 => x"802e8a38",
  1172 => x"870bb6f0",
  1173 => x"0831b6f0",
  1174 => x"0c70b6f8",
  1175 => x"0c738a2a",
  1176 => x"70810651",
  1177 => x"5170802e",
  1178 => x"9238b6ec",
  1179 => x"0851ff71",
  1180 => x"25893870",
  1181 => x"e40cff0b",
  1182 => x"b6ec0c80",
  1183 => x"0bbcdc0c",
  1184 => x"a7ce2da7",
  1185 => x"d52d0290",
  1186 => x"050d0402",
  1187 => x"fc050db6",
  1188 => x"ec085170",
  1189 => x"8024fc38",
  1190 => x"72b6ec0c",
  1191 => x"0284050d",
  1192 => x"0402fc05",
  1193 => x"0da7db2d",
  1194 => x"810bbcdc",
  1195 => x"0ca7d52d",
  1196 => x"bcdc0851",
  1197 => x"70fa3802",
  1198 => x"84050d04",
  1199 => x"02fc050d",
  1200 => x"bca851a2",
  1201 => x"942da2eb",
  1202 => x"51a7ca2d",
  1203 => x"a6f42d81",
  1204 => x"f451a58b",
  1205 => x"2d028405",
  1206 => x"0d0402f4",
  1207 => x"050da6dc",
  1208 => x"04b7c808",
  1209 => x"81f02e09",
  1210 => x"81068938",
  1211 => x"810bb7bc",
  1212 => x"0ca6dc04",
  1213 => x"b7c80881",
  1214 => x"e02e0981",
  1215 => x"06893881",
  1216 => x"0bb7c00c",
  1217 => x"a6dc04b7",
  1218 => x"c80852b7",
  1219 => x"c008802e",
  1220 => x"8838b7c8",
  1221 => x"08818005",
  1222 => x"5271842c",
  1223 => x"728f0653",
  1224 => x"53b7bc08",
  1225 => x"802e9938",
  1226 => x"728429b6",
  1227 => x"fc057213",
  1228 => x"81712b70",
  1229 => x"09730806",
  1230 => x"730c5153",
  1231 => x"53a6d204",
  1232 => x"728429b6",
  1233 => x"fc057213",
  1234 => x"83712b72",
  1235 => x"0807720c",
  1236 => x"5353800b",
  1237 => x"b7c00c80",
  1238 => x"0bb7bc0c",
  1239 => x"bca851a2",
  1240 => x"a72db7c8",
  1241 => x"08ff24fe",
  1242 => x"f838800b",
  1243 => x"b7c80c02",
  1244 => x"8c050d04",
  1245 => x"02f8050d",
  1246 => x"b6fc528f",
  1247 => x"51807270",
  1248 => x"8405540c",
  1249 => x"ff115170",
  1250 => x"8025f238",
  1251 => x"0288050d",
  1252 => x"0402f005",
  1253 => x"0d7551a7",
  1254 => x"db2d7082",
  1255 => x"2cfc06b6",
  1256 => x"fc117210",
  1257 => x"9e067108",
  1258 => x"70722a70",
  1259 => x"83068274",
  1260 => x"2b700974",
  1261 => x"06760c54",
  1262 => x"51565753",
  1263 => x"5153a7d5",
  1264 => x"2d71b7c8",
  1265 => x"0c029005",
  1266 => x"0d047198",
  1267 => x"0c04ffb0",
  1268 => x"08b7c80c",
  1269 => x"04810bff",
  1270 => x"b00c0480",
  1271 => x"0bffb00c",
  1272 => x"0402fc05",
  1273 => x"0d800bb7",
  1274 => x"c40c8051",
  1275 => x"84e52d02",
  1276 => x"84050d04",
  1277 => x"02ec050d",
  1278 => x"76548052",
  1279 => x"870b8815",
  1280 => x"80f52d56",
  1281 => x"53747224",
  1282 => x"8338a053",
  1283 => x"725182ee",
  1284 => x"2d81128b",
  1285 => x"1580f52d",
  1286 => x"54527272",
  1287 => x"25de3802",
  1288 => x"94050d04",
  1289 => x"02f0050d",
  1290 => x"bcf40854",
  1291 => x"81f72d80",
  1292 => x"0bbcf80c",
  1293 => x"7308802e",
  1294 => x"81803882",
  1295 => x"0bb7dc0c",
  1296 => x"bcf8088f",
  1297 => x"06b7d80c",
  1298 => x"73085271",
  1299 => x"832e9638",
  1300 => x"71832689",
  1301 => x"3871812e",
  1302 => x"af38a9a5",
  1303 => x"0471852e",
  1304 => x"9f38a9a5",
  1305 => x"04881480",
  1306 => x"f52d8415",
  1307 => x"08b49853",
  1308 => x"545285f3",
  1309 => x"2d718429",
  1310 => x"13700852",
  1311 => x"52a9a904",
  1312 => x"7351a7f4",
  1313 => x"2da9a504",
  1314 => x"bcf00888",
  1315 => x"15082c70",
  1316 => x"81065152",
  1317 => x"71802e87",
  1318 => x"38b49c51",
  1319 => x"a9a204b4",
  1320 => x"a05185f3",
  1321 => x"2d841408",
  1322 => x"5185f32d",
  1323 => x"bcf80881",
  1324 => x"05bcf80c",
  1325 => x"8c1454a8",
  1326 => x"b4040290",
  1327 => x"050d0471",
  1328 => x"bcf40ca8",
  1329 => x"a42dbcf8",
  1330 => x"08ff05bc",
  1331 => x"fc0c0402",
  1332 => x"ec050dbc",
  1333 => x"f4085580",
  1334 => x"f851a791",
  1335 => x"2db7c808",
  1336 => x"812a7081",
  1337 => x"06515271",
  1338 => x"9b388751",
  1339 => x"a7912db7",
  1340 => x"c808812a",
  1341 => x"70810651",
  1342 => x"5271802e",
  1343 => x"b138aa84",
  1344 => x"04a5da2d",
  1345 => x"8751a791",
  1346 => x"2db7c808",
  1347 => x"f438aa94",
  1348 => x"04a5da2d",
  1349 => x"80f851a7",
  1350 => x"912db7c8",
  1351 => x"08f338b7",
  1352 => x"c4088132",
  1353 => x"70b7c40c",
  1354 => x"70525284",
  1355 => x"e52db7c4",
  1356 => x"08a23880",
  1357 => x"da51a791",
  1358 => x"2d81f551",
  1359 => x"a7912d81",
  1360 => x"f251a791",
  1361 => x"2d81eb51",
  1362 => x"a7912d81",
  1363 => x"f451a791",
  1364 => x"2dae9804",
  1365 => x"81f551a7",
  1366 => x"912db7c8",
  1367 => x"08812a70",
  1368 => x"81065152",
  1369 => x"71802e8f",
  1370 => x"38bcfc08",
  1371 => x"5271802e",
  1372 => x"8638ff12",
  1373 => x"bcfc0c81",
  1374 => x"f251a791",
  1375 => x"2db7c808",
  1376 => x"812a7081",
  1377 => x"06515271",
  1378 => x"802e9538",
  1379 => x"bcf808ff",
  1380 => x"05bcfc08",
  1381 => x"54527272",
  1382 => x"25863881",
  1383 => x"13bcfc0c",
  1384 => x"bcfc0870",
  1385 => x"53547380",
  1386 => x"2e8a388c",
  1387 => x"15ff1555",
  1388 => x"55aba604",
  1389 => x"820bb7dc",
  1390 => x"0c718f06",
  1391 => x"b7d80c81",
  1392 => x"eb51a791",
  1393 => x"2db7c808",
  1394 => x"812a7081",
  1395 => x"06515271",
  1396 => x"802ead38",
  1397 => x"7408852e",
  1398 => x"098106a4",
  1399 => x"38881580",
  1400 => x"f52dff05",
  1401 => x"52718816",
  1402 => x"81b72d71",
  1403 => x"982b5271",
  1404 => x"80258838",
  1405 => x"800b8816",
  1406 => x"81b72d74",
  1407 => x"51a7f42d",
  1408 => x"81f451a7",
  1409 => x"912db7c8",
  1410 => x"08812a70",
  1411 => x"81065152",
  1412 => x"71802eb3",
  1413 => x"38740885",
  1414 => x"2e098106",
  1415 => x"aa388815",
  1416 => x"80f52d81",
  1417 => x"05527188",
  1418 => x"1681b72d",
  1419 => x"7181ff06",
  1420 => x"8b1680f5",
  1421 => x"2d545272",
  1422 => x"72278738",
  1423 => x"72881681",
  1424 => x"b72d7451",
  1425 => x"a7f42d80",
  1426 => x"da51a791",
  1427 => x"2db7c808",
  1428 => x"812a7081",
  1429 => x"06515271",
  1430 => x"802e80fb",
  1431 => x"38bcf408",
  1432 => x"bcfc0855",
  1433 => x"5373802e",
  1434 => x"8a388c13",
  1435 => x"ff155553",
  1436 => x"ace50472",
  1437 => x"08527182",
  1438 => x"2ea63871",
  1439 => x"82268938",
  1440 => x"71812ea5",
  1441 => x"38add704",
  1442 => x"71832ead",
  1443 => x"3871842e",
  1444 => x"09810680",
  1445 => x"c2388813",
  1446 => x"0851a9bf",
  1447 => x"2dadd704",
  1448 => x"88130852",
  1449 => x"712dadd7",
  1450 => x"04810b88",
  1451 => x"14082bbc",
  1452 => x"f00832bc",
  1453 => x"f00cadd4",
  1454 => x"04881380",
  1455 => x"f52d8105",
  1456 => x"8b1480f5",
  1457 => x"2d535471",
  1458 => x"74248338",
  1459 => x"80547388",
  1460 => x"1481b72d",
  1461 => x"a8a42d80",
  1462 => x"54800bb7",
  1463 => x"dc0c738f",
  1464 => x"06b7d80c",
  1465 => x"a05273bc",
  1466 => x"fc082e09",
  1467 => x"81069838",
  1468 => x"bcf808ff",
  1469 => x"05743270",
  1470 => x"09810570",
  1471 => x"72079f2a",
  1472 => x"91713151",
  1473 => x"51535371",
  1474 => x"5182ee2d",
  1475 => x"8114548e",
  1476 => x"7425c638",
  1477 => x"b7c40852",
  1478 => x"71b7c80c",
  1479 => x"0294050d",
  1480 => x"04000000",
  1481 => x"00ffffff",
  1482 => x"ff00ffff",
  1483 => x"ffff00ff",
  1484 => x"ffffff00",
  1485 => x"52657365",
  1486 => x"74000000",
  1487 => x"53617665",
  1488 => x"20616e64",
  1489 => x"20526573",
  1490 => x"65740000",
  1491 => x"4f707469",
  1492 => x"6f6e7320",
  1493 => x"10000000",
  1494 => x"536f756e",
  1495 => x"64201000",
  1496 => x"54757262",
  1497 => x"6f000000",
  1498 => x"4d6f7573",
  1499 => x"6520656d",
  1500 => x"756c6174",
  1501 => x"696f6e00",
  1502 => x"45786974",
  1503 => x"00000000",
  1504 => x"4d617374",
  1505 => x"65720000",
  1506 => x"4f504c4c",
  1507 => x"00000000",
  1508 => x"53434300",
  1509 => x"50534700",
  1510 => x"4261636b",
  1511 => x"00000000",
  1512 => x"5363616e",
  1513 => x"6c696e65",
  1514 => x"73000000",
  1515 => x"53442043",
  1516 => x"61726400",
  1517 => x"4a617061",
  1518 => x"6e657365",
  1519 => x"206b6579",
  1520 => x"206c6179",
  1521 => x"6f757400",
  1522 => x"32303438",
  1523 => x"4c422052",
  1524 => x"414d0000",
  1525 => x"34303936",
  1526 => x"4b422052",
  1527 => x"414d0000",
  1528 => x"536c323a",
  1529 => x"204e6f6e",
  1530 => x"65000000",
  1531 => x"536c323a",
  1532 => x"20455345",
  1533 => x"2d534343",
  1534 => x"20314d42",
  1535 => x"2f534343",
  1536 => x"2d490000",
  1537 => x"536c323a",
  1538 => x"20455345",
  1539 => x"2d52414d",
  1540 => x"20314d42",
  1541 => x"2f415343",
  1542 => x"49493800",
  1543 => x"536c323a",
  1544 => x"20455345",
  1545 => x"2d52414d",
  1546 => x"20314d42",
  1547 => x"2f415343",
  1548 => x"49493136",
  1549 => x"00000000",
  1550 => x"536c313a",
  1551 => x"204e6f6e",
  1552 => x"65000000",
  1553 => x"536c313a",
  1554 => x"20455345",
  1555 => x"2d534343",
  1556 => x"20314d42",
  1557 => x"2f534343",
  1558 => x"2d490000",
  1559 => x"536c313a",
  1560 => x"204d6567",
  1561 => x"6152414d",
  1562 => x"00000000",
  1563 => x"56474120",
  1564 => x"2d203331",
  1565 => x"4b487a2c",
  1566 => x"20363048",
  1567 => x"7a000000",
  1568 => x"56474120",
  1569 => x"2d203331",
  1570 => x"4b487a2c",
  1571 => x"20353048",
  1572 => x"7a000000",
  1573 => x"5456202d",
  1574 => x"20343830",
  1575 => x"692c2036",
  1576 => x"30487a00",
  1577 => x"496e6974",
  1578 => x"69616c69",
  1579 => x"7a696e67",
  1580 => x"20534420",
  1581 => x"63617264",
  1582 => x"0a000000",
  1583 => x"53444843",
  1584 => x"206e6f74",
  1585 => x"20737570",
  1586 => x"706f7274",
  1587 => x"65643b00",
  1588 => x"46617433",
  1589 => x"32206e6f",
  1590 => x"74207375",
  1591 => x"70706f72",
  1592 => x"7465643b",
  1593 => x"00000000",
  1594 => x"0a646973",
  1595 => x"61626c69",
  1596 => x"6e672053",
  1597 => x"44206361",
  1598 => x"72640a10",
  1599 => x"204f4b0a",
  1600 => x"00000000",
  1601 => x"4f434d53",
  1602 => x"58202020",
  1603 => x"43464700",
  1604 => x"54727969",
  1605 => x"6e67204d",
  1606 => x"53583342",
  1607 => x"494f532e",
  1608 => x"5359530a",
  1609 => x"00000000",
  1610 => x"4d535833",
  1611 => x"42494f53",
  1612 => x"53595300",
  1613 => x"54727969",
  1614 => x"6e672042",
  1615 => x"494f535f",
  1616 => x"4d32502e",
  1617 => x"524f4d0a",
  1618 => x"00000000",
  1619 => x"42494f53",
  1620 => x"5f4d3250",
  1621 => x"524f4d00",
  1622 => x"4c6f6164",
  1623 => x"696e6720",
  1624 => x"42494f53",
  1625 => x"0a000000",
  1626 => x"52656164",
  1627 => x"20666169",
  1628 => x"6c65640a",
  1629 => x"00000000",
  1630 => x"4c6f6164",
  1631 => x"696e6720",
  1632 => x"42494f53",
  1633 => x"20666169",
  1634 => x"6c65640a",
  1635 => x"00000000",
  1636 => x"4d425220",
  1637 => x"6661696c",
  1638 => x"0a000000",
  1639 => x"46415431",
  1640 => x"36202020",
  1641 => x"00000000",
  1642 => x"46415433",
  1643 => x"32202020",
  1644 => x"00000000",
  1645 => x"4e6f2070",
  1646 => x"61727469",
  1647 => x"74696f6e",
  1648 => x"20736967",
  1649 => x"0a000000",
  1650 => x"42616420",
  1651 => x"70617274",
  1652 => x"0a000000",
  1653 => x"53444843",
  1654 => x"20657272",
  1655 => x"6f72210a",
  1656 => x"00000000",
  1657 => x"53442069",
  1658 => x"6e69742e",
  1659 => x"2e2e0a00",
  1660 => x"53442063",
  1661 => x"61726420",
  1662 => x"72657365",
  1663 => x"74206661",
  1664 => x"696c6564",
  1665 => x"210a0000",
  1666 => x"57726974",
  1667 => x"65206661",
  1668 => x"696c6564",
  1669 => x"0a000000",
  1670 => x"16200000",
  1671 => x"14200000",
  1672 => x"15200000",
  1673 => x"00000002",
  1674 => x"00000002",
  1675 => x"00001734",
  1676 => x"0000067f",
  1677 => x"00000002",
  1678 => x"0000173c",
  1679 => x"00000671",
  1680 => x"00000004",
  1681 => x"0000174c",
  1682 => x"00001ad0",
  1683 => x"00000004",
  1684 => x"00001758",
  1685 => x"00001a88",
  1686 => x"00000001",
  1687 => x"00001760",
  1688 => x"00000007",
  1689 => x"00000001",
  1690 => x"00001768",
  1691 => x"0000000a",
  1692 => x"00000002",
  1693 => x"00001778",
  1694 => x"000013e1",
  1695 => x"00000000",
  1696 => x"00000000",
  1697 => x"00000000",
  1698 => x"00000005",
  1699 => x"00001780",
  1700 => x"00000007",
  1701 => x"00000005",
  1702 => x"00001788",
  1703 => x"00000007",
  1704 => x"00000005",
  1705 => x"00001790",
  1706 => x"00000007",
  1707 => x"00000005",
  1708 => x"00001794",
  1709 => x"00000007",
  1710 => x"00000004",
  1711 => x"00001798",
  1712 => x"00001a28",
  1713 => x"00000000",
  1714 => x"00000000",
  1715 => x"00000000",
  1716 => x"00000003",
  1717 => x"00001b60",
  1718 => x"00000003",
  1719 => x"00000001",
  1720 => x"000017a0",
  1721 => x"0000000b",
  1722 => x"00000001",
  1723 => x"000017ac",
  1724 => x"00000002",
  1725 => x"00000003",
  1726 => x"00001b54",
  1727 => x"00000003",
  1728 => x"00000003",
  1729 => x"00001b44",
  1730 => x"00000004",
  1731 => x"00000001",
  1732 => x"000017b4",
  1733 => x"00000006",
  1734 => x"00000003",
  1735 => x"00001b3c",
  1736 => x"00000002",
  1737 => x"00000004",
  1738 => x"00001798",
  1739 => x"00001a28",
  1740 => x"00000000",
  1741 => x"00000000",
  1742 => x"00000000",
  1743 => x"000017c8",
  1744 => x"000017d4",
  1745 => x"000017e0",
  1746 => x"000017ec",
  1747 => x"00001804",
  1748 => x"0000181c",
  1749 => x"00001838",
  1750 => x"00001844",
  1751 => x"0000185c",
  1752 => x"0000186c",
  1753 => x"00001880",
  1754 => x"00001894",
  1755 => x"ffffffff",
  1756 => x"00000003",
  1757 => x"00000000",
  1758 => x"00000000",
  1759 => x"00000000",
  1760 => x"00000000",
  1761 => x"00000000",
  1762 => x"00000000",
  1763 => x"00000000",
  1764 => x"00000000",
  1765 => x"00000000",
  1766 => x"00000000",
  1767 => x"00000000",
  1768 => x"00000000",
  1769 => x"00000000",
  1770 => x"00000000",
  1771 => x"00000000",
  1772 => x"00000000",
  1773 => x"00000000",
  1774 => x"00000000",
  1775 => x"00000000",
  1776 => x"00000000",
  1777 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

