-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"000b0b0b",
     4 => x"0b8c04ff",
     5 => x"0d800404",
     6 => x"00000017",
     7 => x"00000000",
     8 => x"0b0b0bb9",
     9 => x"e0080b0b",
    10 => x"0bb9e408",
    11 => x"0b0b0bb9",
    12 => x"e8080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"b9e80c0b",
    16 => x"0b0bb9e4",
    17 => x"0c0b0b0b",
    18 => x"b9e00c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0bafe4",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"b9e070bf",
    57 => x"98278b38",
    58 => x"80717084",
    59 => x"05530c81",
    60 => x"e2048c51",
    61 => x"8dbd0402",
    62 => x"fc050df8",
    63 => x"80518f0b",
    64 => x"b9f00c9f",
    65 => x"0bb9f40c",
    66 => x"a0717081",
    67 => x"055334b9",
    68 => x"f408ff05",
    69 => x"b9f40cb9",
    70 => x"f4088025",
    71 => x"eb38b9f0",
    72 => x"08ff05b9",
    73 => x"f00cb9f0",
    74 => x"088025d7",
    75 => x"38028405",
    76 => x"0d0402f0",
    77 => x"050df880",
    78 => x"53f8a054",
    79 => x"83bf5273",
    80 => x"70810555",
    81 => x"33517073",
    82 => x"70810555",
    83 => x"34ff1252",
    84 => x"718025eb",
    85 => x"38fbc053",
    86 => x"9f52a073",
    87 => x"70810555",
    88 => x"34ff1252",
    89 => x"718025f2",
    90 => x"38029005",
    91 => x"0d0402f4",
    92 => x"050d7453",
    93 => x"8e0bb9f0",
    94 => x"08258f38",
    95 => x"82b22db9",
    96 => x"f008ff05",
    97 => x"b9f00c82",
    98 => x"f404b9f0",
    99 => x"08b9f408",
   100 => x"5351728a",
   101 => x"2e098106",
   102 => x"b7387151",
   103 => x"719f24a0",
   104 => x"38b9f008",
   105 => x"a02911f8",
   106 => x"80115151",
   107 => x"a07134b9",
   108 => x"f4088105",
   109 => x"b9f40cb9",
   110 => x"f408519f",
   111 => x"7125e238",
   112 => x"800bb9f4",
   113 => x"0cb9f008",
   114 => x"8105b9f0",
   115 => x"0c83e404",
   116 => x"70a02912",
   117 => x"f8801151",
   118 => x"51727134",
   119 => x"b9f40881",
   120 => x"05b9f40c",
   121 => x"b9f408a0",
   122 => x"2e098106",
   123 => x"8e38800b",
   124 => x"b9f40cb9",
   125 => x"f0088105",
   126 => x"b9f00c02",
   127 => x"8c050d04",
   128 => x"02e8050d",
   129 => x"77795656",
   130 => x"880bfc16",
   131 => x"77712c8f",
   132 => x"06545254",
   133 => x"80537272",
   134 => x"25953871",
   135 => x"53fbe014",
   136 => x"51877134",
   137 => x"8114ff14",
   138 => x"545472f1",
   139 => x"387153f9",
   140 => x"1576712c",
   141 => x"87065351",
   142 => x"71802e8b",
   143 => x"38fbe014",
   144 => x"51717134",
   145 => x"81145472",
   146 => x"8e249538",
   147 => x"8f733153",
   148 => x"fbe01451",
   149 => x"a0713481",
   150 => x"14ff1454",
   151 => x"5472f138",
   152 => x"0298050d",
   153 => x"0402ec05",
   154 => x"0d800bb9",
   155 => x"f80cf68c",
   156 => x"08f69008",
   157 => x"71882c56",
   158 => x"5481ff06",
   159 => x"52737225",
   160 => x"88387154",
   161 => x"820bb9f8",
   162 => x"0c72882c",
   163 => x"7381ff06",
   164 => x"54557473",
   165 => x"258b3872",
   166 => x"b9f80884",
   167 => x"07b9f80c",
   168 => x"5573842b",
   169 => x"86a07125",
   170 => x"83713170",
   171 => x"0b0b0bb6",
   172 => x"a40c8171",
   173 => x"2bff05f6",
   174 => x"880cfecc",
   175 => x"13ff122c",
   176 => x"788829ff",
   177 => x"94057081",
   178 => x"2cb9f808",
   179 => x"52585255",
   180 => x"51525476",
   181 => x"802e8538",
   182 => x"70810751",
   183 => x"70f6940c",
   184 => x"71098105",
   185 => x"f6800c72",
   186 => x"098105f6",
   187 => x"840c0294",
   188 => x"050d0402",
   189 => x"f4050d74",
   190 => x"53727081",
   191 => x"055480f5",
   192 => x"2d527180",
   193 => x"2e893871",
   194 => x"5182ee2d",
   195 => x"85f90402",
   196 => x"8c050d04",
   197 => x"02f8050d",
   198 => x"a6fc2d80",
   199 => x"da51a8b3",
   200 => x"2db9e008",
   201 => x"812a7081",
   202 => x"06515271",
   203 => x"802ee938",
   204 => x"0288050d",
   205 => x"0402f405",
   206 => x"0dbf8808",
   207 => x"99c406b8",
   208 => x"bc0b80f5",
   209 => x"2d525270",
   210 => x"802e8638",
   211 => x"71848007",
   212 => x"52b7f40b",
   213 => x"80f52d72",
   214 => x"07b8980b",
   215 => x"80f52d70",
   216 => x"812a7081",
   217 => x"06515354",
   218 => x"5270802e",
   219 => x"86387182",
   220 => x"80075272",
   221 => x"81065170",
   222 => x"802e8538",
   223 => x"71880752",
   224 => x"b8a40b80",
   225 => x"f52d7084",
   226 => x"2b730781",
   227 => x"8432b9e0",
   228 => x"0c51028c",
   229 => x"050d0402",
   230 => x"f4050d74",
   231 => x"70818432",
   232 => x"bf880c70",
   233 => x"83065253",
   234 => x"70b7ec0b",
   235 => x"880581b7",
   236 => x"2d72892a",
   237 => x"70810651",
   238 => x"5170b8bc",
   239 => x"0b81b72d",
   240 => x"72832a81",
   241 => x"0673882a",
   242 => x"70810651",
   243 => x"52527080",
   244 => x"2e853871",
   245 => x"82075271",
   246 => x"b8980b81",
   247 => x"b72d7284",
   248 => x"2c708306",
   249 => x"515170b8",
   250 => x"a40b81b7",
   251 => x"2d70b9e0",
   252 => x"0c028c05",
   253 => x"0d0402f4",
   254 => x"050db7a4",
   255 => x"0b881180",
   256 => x"f52d8c12",
   257 => x"881180f5",
   258 => x"2d70842b",
   259 => x"73078c13",
   260 => x"881180f5",
   261 => x"2d70882b",
   262 => x"73079413",
   263 => x"80f52d70",
   264 => x"8c2b7207",
   265 => x"b9e00c53",
   266 => x"53535353",
   267 => x"56525351",
   268 => x"028c050d",
   269 => x"04b6f80b",
   270 => x"80f52db9",
   271 => x"e00c0402",
   272 => x"f4050d74",
   273 => x"b7a47187",
   274 => x"06555351",
   275 => x"72881381",
   276 => x"b72d8c12",
   277 => x"71842c70",
   278 => x"87065552",
   279 => x"52728813",
   280 => x"81b72d8c",
   281 => x"1271842c",
   282 => x"70870655",
   283 => x"52527288",
   284 => x"1381b72d",
   285 => x"70842c70",
   286 => x"87065151",
   287 => x"70941381",
   288 => x"b72d028c",
   289 => x"050d0402",
   290 => x"fc050d02",
   291 => x"8b0580f5",
   292 => x"2db6f80b",
   293 => x"81b72d70",
   294 => x"b9e00c02",
   295 => x"84050d04",
   296 => x"02d4050d",
   297 => x"7cb3a452",
   298 => x"5585f32d",
   299 => x"9ea42db9",
   300 => x"e008802e",
   301 => x"83ad3886",
   302 => x"b52db9e0",
   303 => x"085390ed",
   304 => x"2db9e008",
   305 => x"54b9e008",
   306 => x"802e8399",
   307 => x"38a2a72d",
   308 => x"b9e00880",
   309 => x"2e8738b3",
   310 => x"bc5189ea",
   311 => x"049a902d",
   312 => x"b9e00880",
   313 => x"2ea238b3",
   314 => x"d05185f3",
   315 => x"2db3e851",
   316 => x"85f32d86",
   317 => x"942d7284",
   318 => x"0753810b",
   319 => x"fec40c72",
   320 => x"fec00c72",
   321 => x"5187972d",
   322 => x"840bfec4",
   323 => x"0cb48452",
   324 => x"ba805196",
   325 => x"ff2db9e0",
   326 => x"08802e80",
   327 => x"ec387482",
   328 => x"2e098106",
   329 => x"b83872ba",
   330 => x"8c0c87f6",
   331 => x"2db9e008",
   332 => x"ba900c88",
   333 => x"b52db9e0",
   334 => x"08ba940c",
   335 => x"ba985480",
   336 => x"fc538074",
   337 => x"70840556",
   338 => x"0cff1353",
   339 => x"728025f2",
   340 => x"38ba8c52",
   341 => x"ba805199",
   342 => x"ea2d8b89",
   343 => x"0474812e",
   344 => x"098106a5",
   345 => x"38ba8c52",
   346 => x"ba805199",
   347 => x"c42dba8c",
   348 => x"08ba9008",
   349 => x"525388bf",
   350 => x"2dba9408",
   351 => x"5189872d",
   352 => x"72fec00c",
   353 => x"72518797",
   354 => x"2db49051",
   355 => x"85f32db4",
   356 => x"a852ba80",
   357 => x"5196ff2d",
   358 => x"b9e00898",
   359 => x"38b4b451",
   360 => x"85f32db4",
   361 => x"cc52ba80",
   362 => x"5196ff2d",
   363 => x"b9e00880",
   364 => x"2e81b038",
   365 => x"b4d85185",
   366 => x"f32dba84",
   367 => x"08578077",
   368 => x"595a767a",
   369 => x"2e8b3881",
   370 => x"1a78812a",
   371 => x"595a77f7",
   372 => x"38f71a5a",
   373 => x"80772581",
   374 => x"80387952",
   375 => x"77518480",
   376 => x"2dba8c52",
   377 => x"ba805199",
   378 => x"c42db9e0",
   379 => x"0853b9e0",
   380 => x"08802e80",
   381 => x"c938ba8c",
   382 => x"5b80598c",
   383 => x"ab047a70",
   384 => x"84055c08",
   385 => x"7081ff06",
   386 => x"71882c70",
   387 => x"81ff0673",
   388 => x"902c7081",
   389 => x"ff067598",
   390 => x"2afec80c",
   391 => x"fec80c58",
   392 => x"fec80c57",
   393 => x"fec80c84",
   394 => x"1a5a5376",
   395 => x"53848077",
   396 => x"25843884",
   397 => x"80537279",
   398 => x"24c4388c",
   399 => x"c904b4e8",
   400 => x"5185f32d",
   401 => x"72548ce5",
   402 => x"04ba8051",
   403 => x"99972dfc",
   404 => x"80178119",
   405 => x"59578bd4",
   406 => x"04820bfe",
   407 => x"c40c8154",
   408 => x"8ce50480",
   409 => x"5473b9e0",
   410 => x"0c02ac05",
   411 => x"0d0402f8",
   412 => x"050da983",
   413 => x"2d81f72d",
   414 => x"815184e5",
   415 => x"2dfec452",
   416 => x"81720ca5",
   417 => x"fc2da5fc",
   418 => x"2d84720c",
   419 => x"735189a0",
   420 => x"2db6a851",
   421 => x"aae12d80",
   422 => x"5184e52d",
   423 => x"0288050d",
   424 => x"0402fc05",
   425 => x"0d82518c",
   426 => x"ee2d0284",
   427 => x"050d0402",
   428 => x"fc050d80",
   429 => x"518cee2d",
   430 => x"0284050d",
   431 => x"0402ec05",
   432 => x"0d84b851",
   433 => x"87972d81",
   434 => x"0bfec40c",
   435 => x"84b80bfe",
   436 => x"c00c840b",
   437 => x"fec40c83",
   438 => x"0bfecc0c",
   439 => x"81eef751",
   440 => x"88bf2d87",
   441 => x"f62db9e0",
   442 => x"08fed40c",
   443 => x"a6972da8",
   444 => x"f72da5fc",
   445 => x"2da5fc2d",
   446 => x"81f72d81",
   447 => x"5184e52d",
   448 => x"a5fc2da5",
   449 => x"fc2d8151",
   450 => x"84e52d81",
   451 => x"5189a02d",
   452 => x"b9e00880",
   453 => x"2e828338",
   454 => x"805184e5",
   455 => x"2db6a851",
   456 => x"aae12dbe",
   457 => x"e8085271",
   458 => x"8b38beec",
   459 => x"08527180",
   460 => x"2e818f38",
   461 => x"fed00870",
   462 => x"81065152",
   463 => x"71802e81",
   464 => x"8138a8fd",
   465 => x"2dbee808",
   466 => x"beec0854",
   467 => x"5480ff74",
   468 => x"25843880",
   469 => x"ff5480ff",
   470 => x"73258438",
   471 => x"80ff5373",
   472 => x"ff802584",
   473 => x"38ff8054",
   474 => x"72ff8025",
   475 => x"8438ff80",
   476 => x"53bee808",
   477 => x"707531be",
   478 => x"e80c52be",
   479 => x"ec087074",
   480 => x"31beec0c",
   481 => x"52a8f72d",
   482 => x"b6f80b80",
   483 => x"f52d7081",
   484 => x"2a708106",
   485 => x"51535571",
   486 => x"802e8938",
   487 => x"73812c73",
   488 => x"812c5454",
   489 => x"74810652",
   490 => x"71802e85",
   491 => x"3872812c",
   492 => x"5373882b",
   493 => x"83fe8006",
   494 => x"7381ff06",
   495 => x"7107fed0",
   496 => x"0c52a6fc",
   497 => x"2daaf12d",
   498 => x"b9e00853",
   499 => x"86b52db9",
   500 => x"e008fec0",
   501 => x"0c87f62d",
   502 => x"b9e008fe",
   503 => x"d40c86b5",
   504 => x"2db9e008",
   505 => x"b9fc082e",
   506 => x"9c38b9e0",
   507 => x"08b9fc0c",
   508 => x"84527251",
   509 => x"84e52da5",
   510 => x"fc2da5fc",
   511 => x"2dff1252",
   512 => x"718025ee",
   513 => x"3872802e",
   514 => x"89388a0b",
   515 => x"fec40c8e",
   516 => x"a304820b",
   517 => x"fec40c8e",
   518 => x"a304b4f8",
   519 => x"5185f32d",
   520 => x"820bfec4",
   521 => x"0c800bb9",
   522 => x"e00c0294",
   523 => x"050d0402",
   524 => x"e8050d77",
   525 => x"797b5855",
   526 => x"55805372",
   527 => x"7625a338",
   528 => x"74708105",
   529 => x"5680f52d",
   530 => x"74708105",
   531 => x"5680f52d",
   532 => x"52527171",
   533 => x"2e863881",
   534 => x"5190e404",
   535 => x"81135390",
   536 => x"bb048051",
   537 => x"70b9e00c",
   538 => x"0298050d",
   539 => x"0402d805",
   540 => x"0d800bbe",
   541 => x"940cba8c",
   542 => x"528051a1",
   543 => x"8c2db9e0",
   544 => x"0854b9e0",
   545 => x"088c38b5",
   546 => x"905185f3",
   547 => x"2d735596",
   548 => x"88048056",
   549 => x"810bbeb8",
   550 => x"0c8853b5",
   551 => x"9c52bac2",
   552 => x"5190af2d",
   553 => x"b9e00876",
   554 => x"2e098106",
   555 => x"8738b9e0",
   556 => x"08beb80c",
   557 => x"8853b5a8",
   558 => x"52bade51",
   559 => x"90af2db9",
   560 => x"e0088738",
   561 => x"b9e008be",
   562 => x"b80cbeb8",
   563 => x"08802e80",
   564 => x"f638bdd2",
   565 => x"0b80f52d",
   566 => x"bdd30b80",
   567 => x"f52d7198",
   568 => x"2b71902b",
   569 => x"07bdd40b",
   570 => x"80f52d70",
   571 => x"882b7207",
   572 => x"bdd50b80",
   573 => x"f52d7107",
   574 => x"be8a0b80",
   575 => x"f52dbe8b",
   576 => x"0b80f52d",
   577 => x"71882b07",
   578 => x"535f5452",
   579 => x"5a565755",
   580 => x"7381abaa",
   581 => x"2e098106",
   582 => x"8d387551",
   583 => x"a2ae2db9",
   584 => x"e0085692",
   585 => x"b3047382",
   586 => x"d4d52e87",
   587 => x"38b5b451",
   588 => x"92f404ba",
   589 => x"8c527551",
   590 => x"a18c2db9",
   591 => x"e00855b9",
   592 => x"e008802e",
   593 => x"83c23888",
   594 => x"53b5a852",
   595 => x"bade5190",
   596 => x"af2db9e0",
   597 => x"08893881",
   598 => x"0bbe940c",
   599 => x"92fa0488",
   600 => x"53b59c52",
   601 => x"bac25190",
   602 => x"af2db9e0",
   603 => x"08802e8a",
   604 => x"38b5c851",
   605 => x"85f32d93",
   606 => x"d404be8a",
   607 => x"0b80f52d",
   608 => x"547380d5",
   609 => x"2e098106",
   610 => x"80ca38be",
   611 => x"8b0b80f5",
   612 => x"2d547381",
   613 => x"aa2e0981",
   614 => x"06ba3880",
   615 => x"0bba8c0b",
   616 => x"80f52d56",
   617 => x"547481e9",
   618 => x"2e833881",
   619 => x"547481eb",
   620 => x"2e8c3880",
   621 => x"5573752e",
   622 => x"09810682",
   623 => x"cb38ba97",
   624 => x"0b80f52d",
   625 => x"55748d38",
   626 => x"ba980b80",
   627 => x"f52d5473",
   628 => x"822e8638",
   629 => x"80559688",
   630 => x"04ba990b",
   631 => x"80f52d70",
   632 => x"be8c0cff",
   633 => x"05be900c",
   634 => x"ba9a0b80",
   635 => x"f52dba9b",
   636 => x"0b80f52d",
   637 => x"58760577",
   638 => x"82802905",
   639 => x"70be980c",
   640 => x"ba9c0b80",
   641 => x"f52d70be",
   642 => x"ac0cbe94",
   643 => x"08595758",
   644 => x"76802e81",
   645 => x"a3388853",
   646 => x"b5a852ba",
   647 => x"de5190af",
   648 => x"2db9e008",
   649 => x"81e238be",
   650 => x"8c087084",
   651 => x"2bbeb00c",
   652 => x"70bea80c",
   653 => x"bab10b80",
   654 => x"f52dbab0",
   655 => x"0b80f52d",
   656 => x"71828029",
   657 => x"05bab20b",
   658 => x"80f52d70",
   659 => x"84808029",
   660 => x"12bab30b",
   661 => x"80f52d70",
   662 => x"81800a29",
   663 => x"1270beb4",
   664 => x"0cbeac08",
   665 => x"7129be98",
   666 => x"080570be",
   667 => x"9c0cbab9",
   668 => x"0b80f52d",
   669 => x"bab80b80",
   670 => x"f52d7182",
   671 => x"802905ba",
   672 => x"ba0b80f5",
   673 => x"2d708480",
   674 => x"802912ba",
   675 => x"bb0b80f5",
   676 => x"2d70982b",
   677 => x"81f00a06",
   678 => x"720570be",
   679 => x"a00cfe11",
   680 => x"7e297705",
   681 => x"bea40c52",
   682 => x"59524354",
   683 => x"5e515259",
   684 => x"525d5759",
   685 => x"57968604",
   686 => x"ba9e0b80",
   687 => x"f52dba9d",
   688 => x"0b80f52d",
   689 => x"71828029",
   690 => x"0570beb0",
   691 => x"0c70a029",
   692 => x"83ff0570",
   693 => x"892a70be",
   694 => x"a80cbaa3",
   695 => x"0b80f52d",
   696 => x"baa20b80",
   697 => x"f52d7182",
   698 => x"80290570",
   699 => x"beb40c7b",
   700 => x"71291e70",
   701 => x"bea40c7d",
   702 => x"bea00c73",
   703 => x"05be9c0c",
   704 => x"555e5151",
   705 => x"55558155",
   706 => x"74b9e00c",
   707 => x"02a8050d",
   708 => x"0402ec05",
   709 => x"0d767087",
   710 => x"2c7180ff",
   711 => x"06555654",
   712 => x"be94088a",
   713 => x"3873882c",
   714 => x"7481ff06",
   715 => x"5455ba8c",
   716 => x"52be9808",
   717 => x"1551a18c",
   718 => x"2db9e008",
   719 => x"54b9e008",
   720 => x"802eb338",
   721 => x"be940880",
   722 => x"2e983872",
   723 => x"8429ba8c",
   724 => x"05700852",
   725 => x"53a2ae2d",
   726 => x"b9e008f0",
   727 => x"0a065396",
   728 => x"f4047210",
   729 => x"ba8c0570",
   730 => x"80e02d52",
   731 => x"53a2de2d",
   732 => x"b9e00853",
   733 => x"725473b9",
   734 => x"e00c0294",
   735 => x"050d0402",
   736 => x"c8050d7f",
   737 => x"615f5b80",
   738 => x"0bbea008",
   739 => x"bea40859",
   740 => x"5d56be94",
   741 => x"08762e8a",
   742 => x"38be8c08",
   743 => x"842b5897",
   744 => x"a804bea8",
   745 => x"08842b58",
   746 => x"80597878",
   747 => x"2781a938",
   748 => x"788f06a0",
   749 => x"17575473",
   750 => x"8f38ba8c",
   751 => x"52765181",
   752 => x"1757a18c",
   753 => x"2dba8c56",
   754 => x"807680f5",
   755 => x"2d565474",
   756 => x"742e8338",
   757 => x"81547481",
   758 => x"e52e80f6",
   759 => x"38817075",
   760 => x"06555d73",
   761 => x"802e80ea",
   762 => x"388b1680",
   763 => x"f52d9806",
   764 => x"5a7980de",
   765 => x"388b537d",
   766 => x"52755190",
   767 => x"af2db9e0",
   768 => x"0880cf38",
   769 => x"9c160851",
   770 => x"a2ae2db9",
   771 => x"e008841c",
   772 => x"0c9a1680",
   773 => x"e02d51a2",
   774 => x"de2db9e0",
   775 => x"08b9e008",
   776 => x"881d0cb9",
   777 => x"e0085555",
   778 => x"be940880",
   779 => x"2e983894",
   780 => x"1680e02d",
   781 => x"51a2de2d",
   782 => x"b9e00890",
   783 => x"2b83fff0",
   784 => x"0a067016",
   785 => x"51547388",
   786 => x"1c0c797b",
   787 => x"0c7c5499",
   788 => x"8e048119",
   789 => x"5997aa04",
   790 => x"be940880",
   791 => x"2eae387b",
   792 => x"5196912d",
   793 => x"b9e008b9",
   794 => x"e00880ff",
   795 => x"fffff806",
   796 => x"555c7380",
   797 => x"fffffff8",
   798 => x"2e9238b9",
   799 => x"e008fe05",
   800 => x"be8c0829",
   801 => x"be9c0805",
   802 => x"5797a804",
   803 => x"805473b9",
   804 => x"e00c02b8",
   805 => x"050d0402",
   806 => x"f4050d74",
   807 => x"70088105",
   808 => x"710c7008",
   809 => x"be900806",
   810 => x"5353718e",
   811 => x"38881308",
   812 => x"5196912d",
   813 => x"b9e00888",
   814 => x"140c810b",
   815 => x"b9e00c02",
   816 => x"8c050d04",
   817 => x"02f0050d",
   818 => x"75881108",
   819 => x"fe05be8c",
   820 => x"0829be9c",
   821 => x"08117208",
   822 => x"be900806",
   823 => x"05795553",
   824 => x"5454a18c",
   825 => x"2d029005",
   826 => x"0d0402f0",
   827 => x"050d7588",
   828 => x"1108fe05",
   829 => x"be8c0829",
   830 => x"be9c0811",
   831 => x"7208be90",
   832 => x"08060579",
   833 => x"55535454",
   834 => x"9fcc2d02",
   835 => x"90050d04",
   836 => x"be9408b9",
   837 => x"e00c0402",
   838 => x"f4050dd4",
   839 => x"5281ff72",
   840 => x"0c710853",
   841 => x"81ff720c",
   842 => x"72882b83",
   843 => x"fe800672",
   844 => x"087081ff",
   845 => x"06515253",
   846 => x"81ff720c",
   847 => x"72710788",
   848 => x"2b720870",
   849 => x"81ff0651",
   850 => x"525381ff",
   851 => x"720c7271",
   852 => x"07882b72",
   853 => x"087081ff",
   854 => x"067207b9",
   855 => x"e00c5253",
   856 => x"028c050d",
   857 => x"0402f405",
   858 => x"0d747671",
   859 => x"81ff06d4",
   860 => x"0c5353be",
   861 => x"bc088538",
   862 => x"71892b52",
   863 => x"71982ad4",
   864 => x"0c71902a",
   865 => x"7081ff06",
   866 => x"d40c5171",
   867 => x"882a7081",
   868 => x"ff06d40c",
   869 => x"517181ff",
   870 => x"06d40c72",
   871 => x"902a7081",
   872 => x"ff06d40c",
   873 => x"51d40870",
   874 => x"81ff0651",
   875 => x"5182b8bf",
   876 => x"527081ff",
   877 => x"2e098106",
   878 => x"943881ff",
   879 => x"0bd40cd4",
   880 => x"087081ff",
   881 => x"06ff1454",
   882 => x"515171e5",
   883 => x"3870b9e0",
   884 => x"0c028c05",
   885 => x"0d0402fc",
   886 => x"050d81c7",
   887 => x"5181ff0b",
   888 => x"d40cff11",
   889 => x"51708025",
   890 => x"f4380284",
   891 => x"050d0402",
   892 => x"f0050d9b",
   893 => x"d62d8fcf",
   894 => x"53805287",
   895 => x"fc80f751",
   896 => x"9ae52db9",
   897 => x"e00854b9",
   898 => x"e008812e",
   899 => x"098106a3",
   900 => x"3881ff0b",
   901 => x"d40c820a",
   902 => x"52849c80",
   903 => x"e9519ae5",
   904 => x"2db9e008",
   905 => x"8b3881ff",
   906 => x"0bd40c73",
   907 => x"539cb904",
   908 => x"9bd62dff",
   909 => x"135372c1",
   910 => x"3872b9e0",
   911 => x"0c029005",
   912 => x"0d0402f4",
   913 => x"050d81ff",
   914 => x"0bd40c93",
   915 => x"53805287",
   916 => x"fc80c151",
   917 => x"9ae52db9",
   918 => x"e0088b38",
   919 => x"81ff0bd4",
   920 => x"0c81539c",
   921 => x"ef049bd6",
   922 => x"2dff1353",
   923 => x"72df3872",
   924 => x"b9e00c02",
   925 => x"8c050d04",
   926 => x"02f0050d",
   927 => x"9bd62d83",
   928 => x"aa52849c",
   929 => x"80c8519a",
   930 => x"e52db9e0",
   931 => x"08812e09",
   932 => x"81069238",
   933 => x"9a972db9",
   934 => x"e00883ff",
   935 => x"ff065372",
   936 => x"83aa2e97",
   937 => x"389cc22d",
   938 => x"9db60481",
   939 => x"549e9b04",
   940 => x"b5d45185",
   941 => x"f32d8054",
   942 => x"9e9b0481",
   943 => x"ff0bd40c",
   944 => x"b1539bef",
   945 => x"2db9e008",
   946 => x"802e80c0",
   947 => x"38805287",
   948 => x"fc80fa51",
   949 => x"9ae52db9",
   950 => x"e008b138",
   951 => x"81ff0bd4",
   952 => x"0cd40853",
   953 => x"81ff0bd4",
   954 => x"0c81ff0b",
   955 => x"d40c81ff",
   956 => x"0bd40c81",
   957 => x"ff0bd40c",
   958 => x"72862a70",
   959 => x"8106b9e0",
   960 => x"08565153",
   961 => x"72802e93",
   962 => x"389dab04",
   963 => x"72822eff",
   964 => x"9f38ff13",
   965 => x"5372ffaa",
   966 => x"38725473",
   967 => x"b9e00c02",
   968 => x"90050d04",
   969 => x"02f0050d",
   970 => x"810bbebc",
   971 => x"0c8454d0",
   972 => x"08708f2a",
   973 => x"70810651",
   974 => x"515372f3",
   975 => x"3872d00c",
   976 => x"9bd62db5",
   977 => x"e45185f3",
   978 => x"2dd00870",
   979 => x"8f2a7081",
   980 => x"06515153",
   981 => x"72f33881",
   982 => x"0bd00cb1",
   983 => x"53805284",
   984 => x"d480c051",
   985 => x"9ae52db9",
   986 => x"e008812e",
   987 => x"a1387282",
   988 => x"2e098106",
   989 => x"8c38b5f0",
   990 => x"5185f32d",
   991 => x"80539fc3",
   992 => x"04ff1353",
   993 => x"72d738ff",
   994 => x"145473ff",
   995 => x"a2389cf8",
   996 => x"2db9e008",
   997 => x"bebc0cb9",
   998 => x"e0088b38",
   999 => x"815287fc",
  1000 => x"80d0519a",
  1001 => x"e52d81ff",
  1002 => x"0bd40cd0",
  1003 => x"08708f2a",
  1004 => x"70810651",
  1005 => x"515372f3",
  1006 => x"3872d00c",
  1007 => x"81ff0bd4",
  1008 => x"0c815372",
  1009 => x"b9e00c02",
  1010 => x"90050d04",
  1011 => x"02e8050d",
  1012 => x"785681ff",
  1013 => x"0bd40cd0",
  1014 => x"08708f2a",
  1015 => x"70810651",
  1016 => x"515372f3",
  1017 => x"3882810b",
  1018 => x"d00c81ff",
  1019 => x"0bd40c77",
  1020 => x"5287fc80",
  1021 => x"d8519ae5",
  1022 => x"2db9e008",
  1023 => x"802e8c38",
  1024 => x"b6885185",
  1025 => x"f32d8153",
  1026 => x"a1830481",
  1027 => x"ff0bd40c",
  1028 => x"81fe0bd4",
  1029 => x"0c80ff55",
  1030 => x"75708405",
  1031 => x"57087098",
  1032 => x"2ad40c70",
  1033 => x"902c7081",
  1034 => x"ff06d40c",
  1035 => x"5470882c",
  1036 => x"7081ff06",
  1037 => x"d40c5470",
  1038 => x"81ff06d4",
  1039 => x"0c54ff15",
  1040 => x"55748025",
  1041 => x"d33881ff",
  1042 => x"0bd40c81",
  1043 => x"ff0bd40c",
  1044 => x"81ff0bd4",
  1045 => x"0c868da0",
  1046 => x"5481ff0b",
  1047 => x"d40cd408",
  1048 => x"81ff0655",
  1049 => x"748738ff",
  1050 => x"145473ed",
  1051 => x"3881ff0b",
  1052 => x"d40cd008",
  1053 => x"708f2a70",
  1054 => x"81065151",
  1055 => x"5372f338",
  1056 => x"72d00c72",
  1057 => x"b9e00c02",
  1058 => x"98050d04",
  1059 => x"02e8050d",
  1060 => x"78558056",
  1061 => x"81ff0bd4",
  1062 => x"0cd00870",
  1063 => x"8f2a7081",
  1064 => x"06515153",
  1065 => x"72f33882",
  1066 => x"810bd00c",
  1067 => x"81ff0bd4",
  1068 => x"0c775287",
  1069 => x"fc80d151",
  1070 => x"9ae52d80",
  1071 => x"dbc6df54",
  1072 => x"b9e00880",
  1073 => x"2e8a38b4",
  1074 => x"e85185f3",
  1075 => x"2da29e04",
  1076 => x"81ff0bd4",
  1077 => x"0cd40870",
  1078 => x"81ff0651",
  1079 => x"537281fe",
  1080 => x"2e098106",
  1081 => x"9d3880ff",
  1082 => x"539a972d",
  1083 => x"b9e00875",
  1084 => x"70840557",
  1085 => x"0cff1353",
  1086 => x"728025ed",
  1087 => x"388156a2",
  1088 => x"8804ff14",
  1089 => x"5473c938",
  1090 => x"81ff0bd4",
  1091 => x"0cd00870",
  1092 => x"8f2a7081",
  1093 => x"06515153",
  1094 => x"72f33872",
  1095 => x"d00c75b9",
  1096 => x"e00c0298",
  1097 => x"050d04be",
  1098 => x"bc08b9e0",
  1099 => x"0c0402f4",
  1100 => x"050d7470",
  1101 => x"882a83fe",
  1102 => x"80067072",
  1103 => x"982a0772",
  1104 => x"882b87fc",
  1105 => x"80800673",
  1106 => x"982b81f0",
  1107 => x"0a067173",
  1108 => x"0707b9e0",
  1109 => x"0c565153",
  1110 => x"51028c05",
  1111 => x"0d0402f8",
  1112 => x"050d028e",
  1113 => x"0580f52d",
  1114 => x"74882b07",
  1115 => x"7083ffff",
  1116 => x"06b9e00c",
  1117 => x"51028805",
  1118 => x"0d0402fc",
  1119 => x"050d7251",
  1120 => x"80710c80",
  1121 => x"0b84120c",
  1122 => x"0284050d",
  1123 => x"0402f005",
  1124 => x"0d757008",
  1125 => x"84120853",
  1126 => x"5353ff54",
  1127 => x"71712ea8",
  1128 => x"38a8fd2d",
  1129 => x"84130870",
  1130 => x"84291488",
  1131 => x"11700870",
  1132 => x"81ff0684",
  1133 => x"18088111",
  1134 => x"8706841a",
  1135 => x"0c535155",
  1136 => x"515151a8",
  1137 => x"f72d7154",
  1138 => x"73b9e00c",
  1139 => x"0290050d",
  1140 => x"0402f405",
  1141 => x"0da8fd2d",
  1142 => x"e008e408",
  1143 => x"718b2a70",
  1144 => x"81065153",
  1145 => x"54527080",
  1146 => x"2e9d38be",
  1147 => x"c0087084",
  1148 => x"29bec805",
  1149 => x"7381ff06",
  1150 => x"710c5151",
  1151 => x"bec00881",
  1152 => x"118706be",
  1153 => x"c00c5172",
  1154 => x"8b2a7081",
  1155 => x"06515170",
  1156 => x"802e819b",
  1157 => x"38b99008",
  1158 => x"8429bef4",
  1159 => x"057381ff",
  1160 => x"06710c51",
  1161 => x"b9900881",
  1162 => x"05b9900c",
  1163 => x"850bb98c",
  1164 => x"0cb99008",
  1165 => x"b988082e",
  1166 => x"09810681",
  1167 => x"af38800b",
  1168 => x"b9900cbf",
  1169 => x"840881a4",
  1170 => x"38bef408",
  1171 => x"70097083",
  1172 => x"06fecc0c",
  1173 => x"5270852a",
  1174 => x"70810651",
  1175 => x"52527080",
  1176 => x"2e9038be",
  1177 => x"ec08befc",
  1178 => x"08fe8032",
  1179 => x"115151a4",
  1180 => x"fb04beec",
  1181 => x"08befc08",
  1182 => x"11515170",
  1183 => x"beec0c71",
  1184 => x"842a7081",
  1185 => x"06515170",
  1186 => x"802e9338",
  1187 => x"bee808be",
  1188 => x"f80881ff",
  1189 => x"32118111",
  1190 => x"515151a5",
  1191 => x"a804bee8",
  1192 => x"0870bef8",
  1193 => x"08315151",
  1194 => x"70bee80c",
  1195 => x"a5ec04b9",
  1196 => x"8c08ff05",
  1197 => x"b98c0cb9",
  1198 => x"8c08ff2e",
  1199 => x"098106ac",
  1200 => x"38b99008",
  1201 => x"802e9238",
  1202 => x"810bbf84",
  1203 => x"0c870bb9",
  1204 => x"880831b9",
  1205 => x"880ca5e7",
  1206 => x"04bf8408",
  1207 => x"5170802e",
  1208 => x"8638ff11",
  1209 => x"bf840c80",
  1210 => x"0bb9900c",
  1211 => x"800bbef0",
  1212 => x"0ca8f02d",
  1213 => x"a8f72d02",
  1214 => x"8c050d04",
  1215 => x"02fc050d",
  1216 => x"a8fd2d81",
  1217 => x"0bbef00c",
  1218 => x"a8f72dbe",
  1219 => x"f0085170",
  1220 => x"fa380284",
  1221 => x"050d0402",
  1222 => x"f8050dbe",
  1223 => x"c051a2fa",
  1224 => x"2d800bbf",
  1225 => x"840c830b",
  1226 => x"b9880ce4",
  1227 => x"08708c2a",
  1228 => x"70810651",
  1229 => x"51527180",
  1230 => x"2e863884",
  1231 => x"0bb9880c",
  1232 => x"e408708d",
  1233 => x"2a708106",
  1234 => x"51515271",
  1235 => x"802e9f38",
  1236 => x"870bb988",
  1237 => x"0831b988",
  1238 => x"0ce40870",
  1239 => x"8a2a7081",
  1240 => x"06515152",
  1241 => x"71802ef1",
  1242 => x"3881f40b",
  1243 => x"e40ca3d1",
  1244 => x"51a8ec2d",
  1245 => x"a8962d02",
  1246 => x"88050d04",
  1247 => x"02f4050d",
  1248 => x"a7fe04b9",
  1249 => x"e00881f0",
  1250 => x"2e098106",
  1251 => x"8938810b",
  1252 => x"b9d40ca7",
  1253 => x"fe04b9e0",
  1254 => x"0881e02e",
  1255 => x"09810689",
  1256 => x"38810bb9",
  1257 => x"d80ca7fe",
  1258 => x"04b9e008",
  1259 => x"52b9d808",
  1260 => x"802e8838",
  1261 => x"b9e00881",
  1262 => x"80055271",
  1263 => x"842c728f",
  1264 => x"065353b9",
  1265 => x"d408802e",
  1266 => x"99387284",
  1267 => x"29b99405",
  1268 => x"72138171",
  1269 => x"2b700973",
  1270 => x"0806730c",
  1271 => x"515353a7",
  1272 => x"f4047284",
  1273 => x"29b99405",
  1274 => x"72138371",
  1275 => x"2b720807",
  1276 => x"720c5353",
  1277 => x"800bb9d8",
  1278 => x"0c800bb9",
  1279 => x"d40cbec0",
  1280 => x"51a38d2d",
  1281 => x"b9e008ff",
  1282 => x"24fef838",
  1283 => x"800bb9e0",
  1284 => x"0c028c05",
  1285 => x"0d0402f8",
  1286 => x"050db994",
  1287 => x"528f5180",
  1288 => x"72708405",
  1289 => x"540cff11",
  1290 => x"51708025",
  1291 => x"f2380288",
  1292 => x"050d0402",
  1293 => x"f0050d75",
  1294 => x"51a8fd2d",
  1295 => x"70822cfc",
  1296 => x"06b99411",
  1297 => x"72109e06",
  1298 => x"71087072",
  1299 => x"2a708306",
  1300 => x"82742b70",
  1301 => x"09740676",
  1302 => x"0c545156",
  1303 => x"57535153",
  1304 => x"a8f72d71",
  1305 => x"b9e00c02",
  1306 => x"90050d04",
  1307 => x"71980c04",
  1308 => x"ffb008b9",
  1309 => x"e00c0481",
  1310 => x"0bffb00c",
  1311 => x"04800bff",
  1312 => x"b00c0402",
  1313 => x"fc050d80",
  1314 => x"0bb9dc0c",
  1315 => x"805184e5",
  1316 => x"2d028405",
  1317 => x"0d0402ec",
  1318 => x"050d7654",
  1319 => x"8052870b",
  1320 => x"881580f5",
  1321 => x"2d565374",
  1322 => x"72248338",
  1323 => x"a0537251",
  1324 => x"82ee2d81",
  1325 => x"128b1580",
  1326 => x"f52d5452",
  1327 => x"727225de",
  1328 => x"38029405",
  1329 => x"0d0402f0",
  1330 => x"050dbf8c",
  1331 => x"085481f7",
  1332 => x"2d800bbf",
  1333 => x"900c7308",
  1334 => x"802e8180",
  1335 => x"38820bb9",
  1336 => x"f40cbf90",
  1337 => x"088f06b9",
  1338 => x"f00c7308",
  1339 => x"5271832e",
  1340 => x"96387183",
  1341 => x"26893871",
  1342 => x"812eaf38",
  1343 => x"aac70471",
  1344 => x"852e9f38",
  1345 => x"aac70488",
  1346 => x"1480f52d",
  1347 => x"841508b6",
  1348 => x"98535452",
  1349 => x"85f32d71",
  1350 => x"84291370",
  1351 => x"085252aa",
  1352 => x"cb047351",
  1353 => x"a9962daa",
  1354 => x"c704bf88",
  1355 => x"08881508",
  1356 => x"2c708106",
  1357 => x"51527180",
  1358 => x"2e8738b6",
  1359 => x"9c51aac4",
  1360 => x"04b6a051",
  1361 => x"85f32d84",
  1362 => x"14085185",
  1363 => x"f32dbf90",
  1364 => x"088105bf",
  1365 => x"900c8c14",
  1366 => x"54a9d604",
  1367 => x"0290050d",
  1368 => x"0471bf8c",
  1369 => x"0ca9c62d",
  1370 => x"bf9008ff",
  1371 => x"05bf940c",
  1372 => x"0402e805",
  1373 => x"0d800bbf",
  1374 => x"8c085656",
  1375 => x"80f851a8",
  1376 => x"b32db9e0",
  1377 => x"08812a70",
  1378 => x"81065152",
  1379 => x"71762e09",
  1380 => x"81069b38",
  1381 => x"8751a8b3",
  1382 => x"2db9e008",
  1383 => x"812a7081",
  1384 => x"06515271",
  1385 => x"762eba38",
  1386 => x"abae04a6",
  1387 => x"fc2d8751",
  1388 => x"a8b32db9",
  1389 => x"e008f438",
  1390 => x"abbe04a6",
  1391 => x"fc2d80f8",
  1392 => x"51a8b32d",
  1393 => x"b9e008f3",
  1394 => x"38b9dc08",
  1395 => x"813270b9",
  1396 => x"dc0c7052",
  1397 => x"5284e52d",
  1398 => x"b9dc0880",
  1399 => x"2e833881",
  1400 => x"56b9dc08",
  1401 => x"a23880da",
  1402 => x"51a8b32d",
  1403 => x"81f551a8",
  1404 => x"b32d81f2",
  1405 => x"51a8b32d",
  1406 => x"81eb51a8",
  1407 => x"b32d81f4",
  1408 => x"51a8b32d",
  1409 => x"afdb0481",
  1410 => x"f551a8b3",
  1411 => x"2db9e008",
  1412 => x"812a7081",
  1413 => x"06515271",
  1414 => x"802e9138",
  1415 => x"bf940852",
  1416 => x"71802e88",
  1417 => x"38ff12bf",
  1418 => x"940c8156",
  1419 => x"81f251a8",
  1420 => x"b32db9e0",
  1421 => x"08812a70",
  1422 => x"81065152",
  1423 => x"71802e97",
  1424 => x"38bf9008",
  1425 => x"ff05bf94",
  1426 => x"08545272",
  1427 => x"72258838",
  1428 => x"8113bf94",
  1429 => x"0c8156bf",
  1430 => x"94087053",
  1431 => x"5473802e",
  1432 => x"8a388c15",
  1433 => x"ff155555",
  1434 => x"acdd0482",
  1435 => x"0bb9f40c",
  1436 => x"718f06b9",
  1437 => x"f00c81eb",
  1438 => x"51a8b32d",
  1439 => x"b9e00881",
  1440 => x"2a708106",
  1441 => x"51527180",
  1442 => x"2eaf3881",
  1443 => x"56740885",
  1444 => x"2e098106",
  1445 => x"a4388815",
  1446 => x"80f52dff",
  1447 => x"05527188",
  1448 => x"1681b72d",
  1449 => x"71982b52",
  1450 => x"71802588",
  1451 => x"38800b88",
  1452 => x"1681b72d",
  1453 => x"7451a996",
  1454 => x"2d81f451",
  1455 => x"a8b32db9",
  1456 => x"e008812a",
  1457 => x"70810651",
  1458 => x"5271802e",
  1459 => x"b5388156",
  1460 => x"7408852e",
  1461 => x"098106aa",
  1462 => x"38881580",
  1463 => x"f52d7605",
  1464 => x"52718816",
  1465 => x"81b72d71",
  1466 => x"81ff068b",
  1467 => x"1680f52d",
  1468 => x"54527272",
  1469 => x"27873872",
  1470 => x"881681b7",
  1471 => x"2d7451a9",
  1472 => x"962d80da",
  1473 => x"51a8b32d",
  1474 => x"b9e00881",
  1475 => x"2a708106",
  1476 => x"51527180",
  1477 => x"2e80fe38",
  1478 => x"bf8c08bf",
  1479 => x"94085553",
  1480 => x"73802e8a",
  1481 => x"388c13ff",
  1482 => x"155553ae",
  1483 => x"a0047208",
  1484 => x"5271822e",
  1485 => x"a6387182",
  1486 => x"26893871",
  1487 => x"812ea538",
  1488 => x"af9a0471",
  1489 => x"832ead38",
  1490 => x"71842e09",
  1491 => x"810680ca",
  1492 => x"38881308",
  1493 => x"51aae12d",
  1494 => x"af9a0488",
  1495 => x"13085271",
  1496 => x"2daf9a04",
  1497 => x"810b8814",
  1498 => x"082bbf88",
  1499 => x"0832bf88",
  1500 => x"0caf8f04",
  1501 => x"881380f5",
  1502 => x"2d81058b",
  1503 => x"1480f52d",
  1504 => x"53547174",
  1505 => x"24833880",
  1506 => x"54738814",
  1507 => x"81b72da9",
  1508 => x"c62daf9a",
  1509 => x"0475802e",
  1510 => x"be388054",
  1511 => x"800bb9f4",
  1512 => x"0c738f06",
  1513 => x"b9f00ca0",
  1514 => x"5273bf94",
  1515 => x"082e0981",
  1516 => x"069838bf",
  1517 => x"9008ff05",
  1518 => x"74327009",
  1519 => x"81057072",
  1520 => x"079f2a91",
  1521 => x"71315151",
  1522 => x"53537151",
  1523 => x"82ee2d81",
  1524 => x"14548e74",
  1525 => x"25c638b9",
  1526 => x"dc085271",
  1527 => x"b9e00c02",
  1528 => x"98050d04",
  1529 => x"00ffffff",
  1530 => x"ff00ffff",
  1531 => x"ffff00ff",
  1532 => x"ffffff00",
  1533 => x"52657365",
  1534 => x"74000000",
  1535 => x"53617665",
  1536 => x"20616e64",
  1537 => x"20526573",
  1538 => x"65740000",
  1539 => x"4f707469",
  1540 => x"6f6e7320",
  1541 => x"10000000",
  1542 => x"536f756e",
  1543 => x"64201000",
  1544 => x"54757262",
  1545 => x"6f000000",
  1546 => x"4d6f7573",
  1547 => x"6520456d",
  1548 => x"756c6174",
  1549 => x"696f6e00",
  1550 => x"45786974",
  1551 => x"00000000",
  1552 => x"20205363",
  1553 => x"616c696e",
  1554 => x"6720313a",
  1555 => x"31000000",
  1556 => x"20205363",
  1557 => x"616c696e",
  1558 => x"6720323a",
  1559 => x"31000000",
  1560 => x"20205363",
  1561 => x"616c696e",
  1562 => x"6720323a",
  1563 => x"32000000",
  1564 => x"20205363",
  1565 => x"616c696e",
  1566 => x"6720343a",
  1567 => x"32000000",
  1568 => x"4d617374",
  1569 => x"65720000",
  1570 => x"4f504c4c",
  1571 => x"00000000",
  1572 => x"53434300",
  1573 => x"50534700",
  1574 => x"4261636b",
  1575 => x"00000000",
  1576 => x"5363616e",
  1577 => x"6c696e65",
  1578 => x"73000000",
  1579 => x"53442043",
  1580 => x"61726400",
  1581 => x"4a617061",
  1582 => x"6e657365",
  1583 => x"206b6579",
  1584 => x"206c6179",
  1585 => x"6f757400",
  1586 => x"32303438",
  1587 => x"4b422052",
  1588 => x"414d0000",
  1589 => x"34303936",
  1590 => x"4b422052",
  1591 => x"414d0000",
  1592 => x"536c323a",
  1593 => x"204e6f6e",
  1594 => x"65000000",
  1595 => x"536c323a",
  1596 => x"20455345",
  1597 => x"2d52414d",
  1598 => x"20314d42",
  1599 => x"2f415343",
  1600 => x"49493800",
  1601 => x"536c323a",
  1602 => x"20455345",
  1603 => x"2d534343",
  1604 => x"20314d42",
  1605 => x"2f534343",
  1606 => x"2d490000",
  1607 => x"536c323a",
  1608 => x"20455345",
  1609 => x"2d52414d",
  1610 => x"20314d42",
  1611 => x"2f415343",
  1612 => x"49493136",
  1613 => x"00000000",
  1614 => x"536c313a",
  1615 => x"204e6f6e",
  1616 => x"65000000",
  1617 => x"536c313a",
  1618 => x"20455345",
  1619 => x"2d534343",
  1620 => x"20314d42",
  1621 => x"2f534343",
  1622 => x"2d490000",
  1623 => x"536c313a",
  1624 => x"204d6567",
  1625 => x"6152414d",
  1626 => x"00000000",
  1627 => x"56474120",
  1628 => x"2d203331",
  1629 => x"4b487a2c",
  1630 => x"20363048",
  1631 => x"7a000000",
  1632 => x"56474120",
  1633 => x"2d203331",
  1634 => x"4b487a2c",
  1635 => x"20353048",
  1636 => x"7a000000",
  1637 => x"5456202d",
  1638 => x"20343830",
  1639 => x"692c2036",
  1640 => x"30487a00",
  1641 => x"496e6974",
  1642 => x"69616c69",
  1643 => x"7a696e67",
  1644 => x"20534420",
  1645 => x"63617264",
  1646 => x"0a000000",
  1647 => x"53444843",
  1648 => x"206e6f74",
  1649 => x"20737570",
  1650 => x"706f7274",
  1651 => x"65643b00",
  1652 => x"46617433",
  1653 => x"32206e6f",
  1654 => x"74207375",
  1655 => x"70706f72",
  1656 => x"7465643b",
  1657 => x"00000000",
  1658 => x"0a646973",
  1659 => x"61626c69",
  1660 => x"6e672053",
  1661 => x"44206361",
  1662 => x"72640a10",
  1663 => x"204f4b0a",
  1664 => x"00000000",
  1665 => x"4f434d53",
  1666 => x"58202020",
  1667 => x"43464700",
  1668 => x"54727969",
  1669 => x"6e67204d",
  1670 => x"53583342",
  1671 => x"494f532e",
  1672 => x"5359530a",
  1673 => x"00000000",
  1674 => x"4d535833",
  1675 => x"42494f53",
  1676 => x"53595300",
  1677 => x"54727969",
  1678 => x"6e672042",
  1679 => x"494f535f",
  1680 => x"4d32502e",
  1681 => x"524f4d0a",
  1682 => x"00000000",
  1683 => x"42494f53",
  1684 => x"5f4d3250",
  1685 => x"524f4d00",
  1686 => x"4c6f6164",
  1687 => x"696e6720",
  1688 => x"42494f53",
  1689 => x"0a000000",
  1690 => x"52656164",
  1691 => x"20666169",
  1692 => x"6c65640a",
  1693 => x"00000000",
  1694 => x"4c6f6164",
  1695 => x"696e6720",
  1696 => x"42494f53",
  1697 => x"20666169",
  1698 => x"6c65640a",
  1699 => x"00000000",
  1700 => x"4d425220",
  1701 => x"6661696c",
  1702 => x"0a000000",
  1703 => x"46415431",
  1704 => x"36202020",
  1705 => x"00000000",
  1706 => x"46415433",
  1707 => x"32202020",
  1708 => x"00000000",
  1709 => x"4e6f2070",
  1710 => x"61727469",
  1711 => x"74696f6e",
  1712 => x"20736967",
  1713 => x"0a000000",
  1714 => x"42616420",
  1715 => x"70617274",
  1716 => x"0a000000",
  1717 => x"53444843",
  1718 => x"20657272",
  1719 => x"6f72210a",
  1720 => x"00000000",
  1721 => x"53442069",
  1722 => x"6e69742e",
  1723 => x"2e2e0a00",
  1724 => x"53442063",
  1725 => x"61726420",
  1726 => x"72657365",
  1727 => x"74206661",
  1728 => x"696c6564",
  1729 => x"210a0000",
  1730 => x"57726974",
  1731 => x"65206661",
  1732 => x"696c6564",
  1733 => x"0a000000",
  1734 => x"16200000",
  1735 => x"14200000",
  1736 => x"15200000",
  1737 => x"00000002",
  1738 => x"00000002",
  1739 => x"000017f4",
  1740 => x"000006af",
  1741 => x"00000002",
  1742 => x"000017fc",
  1743 => x"000006a1",
  1744 => x"00000004",
  1745 => x"0000180c",
  1746 => x"00001bec",
  1747 => x"00000004",
  1748 => x"00001818",
  1749 => x"00001ba4",
  1750 => x"00000001",
  1751 => x"00001820",
  1752 => x"00000007",
  1753 => x"00000001",
  1754 => x"00001828",
  1755 => x"0000000a",
  1756 => x"00000003",
  1757 => x"00001b94",
  1758 => x"00000004",
  1759 => x"00000002",
  1760 => x"00001838",
  1761 => x"00001483",
  1762 => x"00000000",
  1763 => x"00000000",
  1764 => x"00000000",
  1765 => x"00001840",
  1766 => x"00001850",
  1767 => x"00001860",
  1768 => x"00001870",
  1769 => x"00000005",
  1770 => x"00001880",
  1771 => x"00000007",
  1772 => x"00000005",
  1773 => x"00001888",
  1774 => x"00000007",
  1775 => x"00000005",
  1776 => x"00001890",
  1777 => x"00000007",
  1778 => x"00000005",
  1779 => x"00001894",
  1780 => x"00000007",
  1781 => x"00000004",
  1782 => x"00001898",
  1783 => x"00001b28",
  1784 => x"00000000",
  1785 => x"00000000",
  1786 => x"00000000",
  1787 => x"00000003",
  1788 => x"00001c7c",
  1789 => x"00000003",
  1790 => x"00000001",
  1791 => x"000018a0",
  1792 => x"0000000b",
  1793 => x"00000001",
  1794 => x"000018ac",
  1795 => x"00000002",
  1796 => x"00000003",
  1797 => x"00001c70",
  1798 => x"00000003",
  1799 => x"00000003",
  1800 => x"00001c60",
  1801 => x"00000004",
  1802 => x"00000001",
  1803 => x"000018b4",
  1804 => x"00000006",
  1805 => x"00000003",
  1806 => x"00001c58",
  1807 => x"00000002",
  1808 => x"00000004",
  1809 => x"00001898",
  1810 => x"00001b28",
  1811 => x"00000000",
  1812 => x"00000000",
  1813 => x"00000000",
  1814 => x"000018c8",
  1815 => x"000018d4",
  1816 => x"000018e0",
  1817 => x"000018ec",
  1818 => x"00001904",
  1819 => x"0000191c",
  1820 => x"00001938",
  1821 => x"00001944",
  1822 => x"0000195c",
  1823 => x"0000196c",
  1824 => x"00001980",
  1825 => x"00001994",
  1826 => x"00000003",
  1827 => x"00000000",
  1828 => x"00000000",
  1829 => x"00000000",
  1830 => x"00000000",
  1831 => x"00000000",
  1832 => x"00000000",
  1833 => x"00000000",
  1834 => x"00000000",
  1835 => x"00000000",
  1836 => x"00000000",
  1837 => x"00000000",
  1838 => x"00000000",
  1839 => x"00000000",
  1840 => x"00000000",
  1841 => x"00000000",
  1842 => x"00000000",
  1843 => x"00000000",
  1844 => x"00000000",
  1845 => x"00000000",
  1846 => x"00000000",
  1847 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

