-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b0bb3",
     9 => x"c0080b0b",
    10 => x"0bb3c408",
    11 => x"0b0b0bb3",
    12 => x"c8080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"b3c80c0b",
    16 => x"0b0bb3c4",
    17 => x"0c0b0b0b",
    18 => x"b3c00c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0ba498",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"b3c070ba",
    57 => x"98278b38",
    58 => x"80717084",
    59 => x"05530c81",
    60 => x"e2048c51",
    61 => x"81f70402",
    62 => x"d8050d81",
    63 => x"0bfec40c",
    64 => x"b90bfec0",
    65 => x"0c840bfe",
    66 => x"c40c9f83",
    67 => x"2da2b12d",
    68 => x"a4a85195",
    69 => x"da2d92f6",
    70 => x"2db3c008",
    71 => x"802e81d2",
    72 => x"3884c92d",
    73 => x"a4c052b4",
    74 => x"f8518b9e",
    75 => x"2db3c008",
    76 => x"81ff0653",
    77 => x"729738a4",
    78 => x"cc52b4f8",
    79 => x"518b9e2d",
    80 => x"b3c00881",
    81 => x"ff065372",
    82 => x"802e81a0",
    83 => x"38a4d851",
    84 => x"95da2db4",
    85 => x"fc085780",
    86 => x"59787725",
    87 => x"819438b5",
    88 => x"9052b4f8",
    89 => x"518df52d",
    90 => x"b3c00881",
    91 => x"ff06b590",
    92 => x"5b538058",
    93 => x"72782e09",
    94 => x"8106b138",
    95 => x"83bf0479",
    96 => x"7084055b",
    97 => x"087081ff",
    98 => x"0671882c",
    99 => x"7081ff06",
   100 => x"73902c70",
   101 => x"81ff0675",
   102 => x"982afec8",
   103 => x"0cfec80c",
   104 => x"58fec80c",
   105 => x"57fec80c",
   106 => x"84195953",
   107 => x"76538480",
   108 => x"77258438",
   109 => x"84805372",
   110 => x"7824c438",
   111 => x"83c504a4",
   112 => x"f45195da",
   113 => x"2db4f851",
   114 => x"8dc82dfc",
   115 => x"8017811a",
   116 => x"5a57ae51",
   117 => x"95b82d78",
   118 => x"bf065372",
   119 => x"86388a51",
   120 => x"95b82d76",
   121 => x"8024fef7",
   122 => x"3883f204",
   123 => x"a5885195",
   124 => x"da2d820b",
   125 => x"fec40c9f",
   126 => x"9b2db3c0",
   127 => x"08802ef7",
   128 => x"38b3c008",
   129 => x"5195b82d",
   130 => x"83f70402",
   131 => x"e8050d77",
   132 => x"797b5855",
   133 => x"55805372",
   134 => x"7625a338",
   135 => x"74708105",
   136 => x"5680f52d",
   137 => x"74708105",
   138 => x"5680f52d",
   139 => x"52527171",
   140 => x"2e863881",
   141 => x"5184c004",
   142 => x"81135384",
   143 => x"97048051",
   144 => x"70b3c00c",
   145 => x"0298050d",
   146 => x"0402d805",
   147 => x"0d800bb9",
   148 => x"a80ca5a0",
   149 => x"5195da2d",
   150 => x"b5905280",
   151 => x"5194952d",
   152 => x"b3c00854",
   153 => x"b3c0088c",
   154 => x"38a5b051",
   155 => x"95da2d73",
   156 => x"558a9c04",
   157 => x"a5c45195",
   158 => x"da2d8056",
   159 => x"810bb584",
   160 => x"0c8853a5",
   161 => x"dc52b5c6",
   162 => x"51848b2d",
   163 => x"b3c00876",
   164 => x"2e098106",
   165 => x"8738b3c0",
   166 => x"08b5840c",
   167 => x"8853a5e8",
   168 => x"52b5e251",
   169 => x"848b2db3",
   170 => x"c0088738",
   171 => x"b3c008b5",
   172 => x"840cb584",
   173 => x"0852a5f4",
   174 => x"5197e22d",
   175 => x"b5840880",
   176 => x"2e818738",
   177 => x"b8d60b80",
   178 => x"f52db8d7",
   179 => x"0b80f52d",
   180 => x"71982b71",
   181 => x"902b07b8",
   182 => x"d80b80f5",
   183 => x"2d70882b",
   184 => x"7207b8d9",
   185 => x"0b80f52d",
   186 => x"7107b98e",
   187 => x"0b80f52d",
   188 => x"b98f0b80",
   189 => x"f52d7188",
   190 => x"2b07535f",
   191 => x"54525a56",
   192 => x"57557381",
   193 => x"abaa2e09",
   194 => x"81068d38",
   195 => x"755196a2",
   196 => x"2db3c008",
   197 => x"5686a804",
   198 => x"7382d4d5",
   199 => x"2e8a38a6",
   200 => x"885195da",
   201 => x"2d87dd04",
   202 => x"7552a6a8",
   203 => x"5197e22d",
   204 => x"b5905275",
   205 => x"5194952d",
   206 => x"b3c00855",
   207 => x"b3c00880",
   208 => x"2e83d938",
   209 => x"a6c05195",
   210 => x"da2da6e8",
   211 => x"5197e22d",
   212 => x"8853a5e8",
   213 => x"52b5e251",
   214 => x"848b2db3",
   215 => x"c0088938",
   216 => x"810bb9a8",
   217 => x"0c878304",
   218 => x"8853a5dc",
   219 => x"52b5c651",
   220 => x"848b2db3",
   221 => x"c008802e",
   222 => x"8a38a780",
   223 => x"5197e22d",
   224 => x"87dd04b9",
   225 => x"8e0b80f5",
   226 => x"2d547380",
   227 => x"d52e0981",
   228 => x"0680ca38",
   229 => x"b98f0b80",
   230 => x"f52d5473",
   231 => x"81aa2e09",
   232 => x"8106ba38",
   233 => x"800bb590",
   234 => x"0b80f52d",
   235 => x"56547481",
   236 => x"e92e8338",
   237 => x"81547481",
   238 => x"eb2e8c38",
   239 => x"80557375",
   240 => x"2e098106",
   241 => x"82d638b5",
   242 => x"9b0b80f5",
   243 => x"2d59788d",
   244 => x"38b59c0b",
   245 => x"80f52d54",
   246 => x"73822e86",
   247 => x"3880558a",
   248 => x"9c04b59d",
   249 => x"0b80f52d",
   250 => x"70b9b00c",
   251 => x"ff1170b9",
   252 => x"a40c5452",
   253 => x"a7a05197",
   254 => x"e22db59e",
   255 => x"0b80f52d",
   256 => x"b59f0b80",
   257 => x"f52d5676",
   258 => x"05758280",
   259 => x"290570b9",
   260 => x"980cb5a0",
   261 => x"0b80f52d",
   262 => x"70b9940c",
   263 => x"b9a80859",
   264 => x"57587680",
   265 => x"2e81a538",
   266 => x"8853a5e8",
   267 => x"52b5e251",
   268 => x"848b2d78",
   269 => x"55b3c008",
   270 => x"81e238b9",
   271 => x"b0087084",
   272 => x"2bb9900c",
   273 => x"70b9ac0c",
   274 => x"b5b50b80",
   275 => x"f52db5b4",
   276 => x"0b80f52d",
   277 => x"71828029",
   278 => x"05b5b60b",
   279 => x"80f52d70",
   280 => x"84808029",
   281 => x"12b5b70b",
   282 => x"80f52d70",
   283 => x"81800a29",
   284 => x"1270b588",
   285 => x"0cb99408",
   286 => x"7129b998",
   287 => x"080570b9",
   288 => x"b80cb5bd",
   289 => x"0b80f52d",
   290 => x"b5bc0b80",
   291 => x"f52d7182",
   292 => x"802905b5",
   293 => x"be0b80f5",
   294 => x"2d708480",
   295 => x"802912b5",
   296 => x"bf0b80f5",
   297 => x"2d70982b",
   298 => x"81f00a06",
   299 => x"720570b5",
   300 => x"8c0cfe11",
   301 => x"7e297705",
   302 => x"b9a00c52",
   303 => x"5752575d",
   304 => x"5751525f",
   305 => x"525c5757",
   306 => x"578a9a04",
   307 => x"b5a20b80",
   308 => x"f52db5a1",
   309 => x"0b80f52d",
   310 => x"71828029",
   311 => x"0570b990",
   312 => x"0c70a029",
   313 => x"83ff0570",
   314 => x"892a70b9",
   315 => x"ac0cb5a7",
   316 => x"0b80f52d",
   317 => x"b5a60b80",
   318 => x"f52d7182",
   319 => x"80290570",
   320 => x"b5880c7b",
   321 => x"71291e70",
   322 => x"b9a00c7d",
   323 => x"b58c0c73",
   324 => x"05b9b80c",
   325 => x"555e5151",
   326 => x"55558155",
   327 => x"74b3c00c",
   328 => x"02a8050d",
   329 => x"0402ec05",
   330 => x"0d767087",
   331 => x"2c7180ff",
   332 => x"06575553",
   333 => x"b9a8088a",
   334 => x"3872882c",
   335 => x"7381ff06",
   336 => x"5654b998",
   337 => x"081452a7",
   338 => x"c45197e2",
   339 => x"2db59052",
   340 => x"b9980814",
   341 => x"5194952d",
   342 => x"b3c00853",
   343 => x"b3c00880",
   344 => x"2eb338b9",
   345 => x"a808802e",
   346 => x"98387484",
   347 => x"29b59005",
   348 => x"70085253",
   349 => x"96a22db3",
   350 => x"c008f00a",
   351 => x"06558b93",
   352 => x"047410b5",
   353 => x"90057080",
   354 => x"e02d5253",
   355 => x"96d22db3",
   356 => x"c0085574",
   357 => x"5372b3c0",
   358 => x"0c029405",
   359 => x"0d0402c8",
   360 => x"050d7f61",
   361 => x"5f5c800b",
   362 => x"b58c08b9",
   363 => x"a0085959",
   364 => x"56b9a808",
   365 => x"762e8a38",
   366 => x"b9b00884",
   367 => x"2b598bc7",
   368 => x"04b9ac08",
   369 => x"842b5980",
   370 => x"5a797927",
   371 => x"81b63879",
   372 => x"8f06a017",
   373 => x"57547397",
   374 => x"387652a7",
   375 => x"e45197e2",
   376 => x"2db59052",
   377 => x"76518117",
   378 => x"5794952d",
   379 => x"b5905680",
   380 => x"7680f52d",
   381 => x"56547474",
   382 => x"2e833881",
   383 => x"547481e5",
   384 => x"2e80fb38",
   385 => x"81707506",
   386 => x"555d7380",
   387 => x"2e80ef38",
   388 => x"8b1680f5",
   389 => x"2d98065b",
   390 => x"7a80e338",
   391 => x"755195da",
   392 => x"2d8b537d",
   393 => x"52755184",
   394 => x"8b2db3c0",
   395 => x"0880cf38",
   396 => x"9c160851",
   397 => x"96a22db3",
   398 => x"c008841d",
   399 => x"0c9a1680",
   400 => x"e02d5196",
   401 => x"d22db3c0",
   402 => x"08b3c008",
   403 => x"881e0cb3",
   404 => x"c0085555",
   405 => x"b9a80880",
   406 => x"2e983894",
   407 => x"1680e02d",
   408 => x"5196d22d",
   409 => x"b3c00890",
   410 => x"2b83fff0",
   411 => x"0a067016",
   412 => x"51547388",
   413 => x"1d0c7a7c",
   414 => x"0c7c548d",
   415 => x"bf04811a",
   416 => x"5a8bc904",
   417 => x"b9a80880",
   418 => x"2eb33877",
   419 => x"518aa52d",
   420 => x"b3c008b3",
   421 => x"c00853a8",
   422 => x"84525897",
   423 => x"e22d7780",
   424 => x"fffffff8",
   425 => x"06547380",
   426 => x"fffffff8",
   427 => x"2e8f38fe",
   428 => x"18b9b008",
   429 => x"29b9b808",
   430 => x"05578bc7",
   431 => x"04805473",
   432 => x"b3c00c02",
   433 => x"b8050d04",
   434 => x"02f4050d",
   435 => x"74700881",
   436 => x"05710c70",
   437 => x"08b9a408",
   438 => x"06535371",
   439 => x"8e388813",
   440 => x"08518aa5",
   441 => x"2db3c008",
   442 => x"88140c81",
   443 => x"0bb3c00c",
   444 => x"028c050d",
   445 => x"0402f005",
   446 => x"0d758811",
   447 => x"08fe05b9",
   448 => x"b00829b9",
   449 => x"b8081172",
   450 => x"08b9a408",
   451 => x"06057955",
   452 => x"53545494",
   453 => x"952db3c0",
   454 => x"0853b3c0",
   455 => x"08802e83",
   456 => x"38815372",
   457 => x"b3c00c02",
   458 => x"90050d04",
   459 => x"02f4050d",
   460 => x"d45281ff",
   461 => x"720c7108",
   462 => x"5381ff72",
   463 => x"0c72882b",
   464 => x"83fe8006",
   465 => x"72087081",
   466 => x"ff065152",
   467 => x"5381ff72",
   468 => x"0c727107",
   469 => x"882b7208",
   470 => x"7081ff06",
   471 => x"51525381",
   472 => x"ff720c72",
   473 => x"7107882b",
   474 => x"72087081",
   475 => x"ff067207",
   476 => x"b3c00c52",
   477 => x"53028c05",
   478 => x"0d0402f4",
   479 => x"050d7476",
   480 => x"7181ff06",
   481 => x"d40c5353",
   482 => x"b9bc0885",
   483 => x"3871892b",
   484 => x"5271982a",
   485 => x"d40c7190",
   486 => x"2a7081ff",
   487 => x"06d40c51",
   488 => x"71882a70",
   489 => x"81ff06d4",
   490 => x"0c517181",
   491 => x"ff06d40c",
   492 => x"72902a70",
   493 => x"81ff06d4",
   494 => x"0c51d408",
   495 => x"7081ff06",
   496 => x"515182b8",
   497 => x"bf527081",
   498 => x"ff2e0981",
   499 => x"06943881",
   500 => x"ff0bd40c",
   501 => x"d4087081",
   502 => x"ff06ff14",
   503 => x"54515171",
   504 => x"e53870b3",
   505 => x"c00c028c",
   506 => x"050d0402",
   507 => x"fc050d81",
   508 => x"c75181ff",
   509 => x"0bd40cff",
   510 => x"11517080",
   511 => x"25f43802",
   512 => x"84050d04",
   513 => x"02f0050d",
   514 => x"8feb2d81",
   515 => x"9c9f5380",
   516 => x"5287fc80",
   517 => x"f7518efa",
   518 => x"2db3c008",
   519 => x"54b3c008",
   520 => x"812e0981",
   521 => x"06a33881",
   522 => x"ff0bd40c",
   523 => x"820a5284",
   524 => x"9c80e951",
   525 => x"8efa2db3",
   526 => x"c0088b38",
   527 => x"81ff0bd4",
   528 => x"0c735390",
   529 => x"cf048feb",
   530 => x"2dff1353",
   531 => x"72c13872",
   532 => x"b3c00c02",
   533 => x"90050d04",
   534 => x"02f4050d",
   535 => x"81ff0bd4",
   536 => x"0ca89c51",
   537 => x"95da2d93",
   538 => x"53805287",
   539 => x"fc80c151",
   540 => x"8efa2db3",
   541 => x"c0088b38",
   542 => x"81ff0bd4",
   543 => x"0c815391",
   544 => x"8b048feb",
   545 => x"2dff1353",
   546 => x"72df3872",
   547 => x"b3c00c02",
   548 => x"8c050d04",
   549 => x"02f0050d",
   550 => x"8feb2d83",
   551 => x"aa52849c",
   552 => x"80c8518e",
   553 => x"fa2db3c0",
   554 => x"08b3c008",
   555 => x"53a8a852",
   556 => x"5397e22d",
   557 => x"72812e09",
   558 => x"81069c38",
   559 => x"8eac2db3",
   560 => x"c00883ff",
   561 => x"ff065372",
   562 => x"83aa2ea1",
   563 => x"38b3c008",
   564 => x"52a8c051",
   565 => x"97e22d90",
   566 => x"d82d91e8",
   567 => x"04815492",
   568 => x"ed04a8d8",
   569 => x"5197e22d",
   570 => x"805492ed",
   571 => x"0481ff0b",
   572 => x"d40cb153",
   573 => x"90842db3",
   574 => x"c008802e",
   575 => x"80e03880",
   576 => x"5287fc80",
   577 => x"fa518efa",
   578 => x"2db3c008",
   579 => x"80c638b3",
   580 => x"c00852a8",
   581 => x"f45197e2",
   582 => x"2d81ff0b",
   583 => x"d40cd408",
   584 => x"7081ff06",
   585 => x"7054a980",
   586 => x"53515397",
   587 => x"e22d81ff",
   588 => x"0bd40c81",
   589 => x"ff0bd40c",
   590 => x"81ff0bd4",
   591 => x"0c81ff0b",
   592 => x"d40c7286",
   593 => x"2a708106",
   594 => x"70565153",
   595 => x"72802e9d",
   596 => x"3891dd04",
   597 => x"b3c00852",
   598 => x"a8f45197",
   599 => x"e22d7282",
   600 => x"2efeff38",
   601 => x"ff135372",
   602 => x"ff8a3872",
   603 => x"5473b3c0",
   604 => x"0c029005",
   605 => x"0d0402f4",
   606 => x"050d810b",
   607 => x"b9bc0cd0",
   608 => x"08708f2a",
   609 => x"70810651",
   610 => x"515372f3",
   611 => x"3872d00c",
   612 => x"8feb2da9",
   613 => x"905195da",
   614 => x"2dd00870",
   615 => x"8f2a7081",
   616 => x"06515153",
   617 => x"72f33881",
   618 => x"0bd00c87",
   619 => x"53805284",
   620 => x"d480c051",
   621 => x"8efa2db3",
   622 => x"c008812e",
   623 => x"94387282",
   624 => x"2e098106",
   625 => x"86388053",
   626 => x"948604ff",
   627 => x"135372dd",
   628 => x"3891942d",
   629 => x"b3c008b9",
   630 => x"bc0cb3c0",
   631 => x"088b3881",
   632 => x"5287fc80",
   633 => x"d0518efa",
   634 => x"2d81ff0b",
   635 => x"d40cd008",
   636 => x"708f2a70",
   637 => x"81065151",
   638 => x"5372f338",
   639 => x"72d00c81",
   640 => x"ff0bd40c",
   641 => x"815372b3",
   642 => x"c00c028c",
   643 => x"050d0480",
   644 => x"0bb3c00c",
   645 => x"0402e005",
   646 => x"0d797b57",
   647 => x"57805881",
   648 => x"ff0bd40c",
   649 => x"d008708f",
   650 => x"2a708106",
   651 => x"51515473",
   652 => x"f3388281",
   653 => x"0bd00c81",
   654 => x"ff0bd40c",
   655 => x"765287fc",
   656 => x"80d1518e",
   657 => x"fa2d80db",
   658 => x"c6df55b3",
   659 => x"c008802e",
   660 => x"9038b3c0",
   661 => x"08537652",
   662 => x"a99c5197",
   663 => x"e22d95af",
   664 => x"0481ff0b",
   665 => x"d40cd408",
   666 => x"7081ff06",
   667 => x"51547381",
   668 => x"fe2e0981",
   669 => x"069d3880",
   670 => x"ff548eac",
   671 => x"2db3c008",
   672 => x"76708405",
   673 => x"580cff14",
   674 => x"54738025",
   675 => x"ed388158",
   676 => x"959904ff",
   677 => x"155574c9",
   678 => x"3881ff0b",
   679 => x"d40cd008",
   680 => x"708f2a70",
   681 => x"81065151",
   682 => x"5473f338",
   683 => x"73d00c77",
   684 => x"b3c00c02",
   685 => x"a0050d04",
   686 => x"02f8050d",
   687 => x"7352c008",
   688 => x"70882a70",
   689 => x"81065151",
   690 => x"5170802e",
   691 => x"f13871c0",
   692 => x"0c71b3c0",
   693 => x"0c028805",
   694 => x"0d0402e8",
   695 => x"050d8078",
   696 => x"57557570",
   697 => x"84055708",
   698 => x"53805472",
   699 => x"982a7388",
   700 => x"2b545271",
   701 => x"802ea238",
   702 => x"c0087088",
   703 => x"2a708106",
   704 => x"51515170",
   705 => x"802ef138",
   706 => x"71c00c81",
   707 => x"15811555",
   708 => x"55837425",
   709 => x"d63871ca",
   710 => x"3874b3c0",
   711 => x"0c029805",
   712 => x"0d0402f4",
   713 => x"050d7470",
   714 => x"882a83fe",
   715 => x"80067072",
   716 => x"982a0772",
   717 => x"882b87fc",
   718 => x"80800673",
   719 => x"982b81f0",
   720 => x"0a067173",
   721 => x"0707b3c0",
   722 => x"0c565153",
   723 => x"51028c05",
   724 => x"0d0402f8",
   725 => x"050d028e",
   726 => x"0580f52d",
   727 => x"74882b07",
   728 => x"7083ffff",
   729 => x"06b3c00c",
   730 => x"51028805",
   731 => x"0d0402f8",
   732 => x"050d7370",
   733 => x"902b7190",
   734 => x"2a07b3c0",
   735 => x"0c520288",
   736 => x"050d0402",
   737 => x"ec050d76",
   738 => x"53805572",
   739 => x"75258b38",
   740 => x"ad5195b8",
   741 => x"2d720981",
   742 => x"05537280",
   743 => x"2eb53887",
   744 => x"54729c2a",
   745 => x"73842b54",
   746 => x"5271802e",
   747 => x"83388155",
   748 => x"89722587",
   749 => x"38b71252",
   750 => x"97be04b0",
   751 => x"12527480",
   752 => x"2e863871",
   753 => x"5195b82d",
   754 => x"ff145473",
   755 => x"8025d238",
   756 => x"97d804b0",
   757 => x"5195b82d",
   758 => x"800bb3c0",
   759 => x"0c029405",
   760 => x"0d0402c0",
   761 => x"050d0280",
   762 => x"c4055780",
   763 => x"70787084",
   764 => x"055a0872",
   765 => x"415f5d58",
   766 => x"7c708405",
   767 => x"5e085a80",
   768 => x"5b79982a",
   769 => x"7a882b5b",
   770 => x"56758638",
   771 => x"775f99da",
   772 => x"047d802e",
   773 => x"81a23880",
   774 => x"5e7580e4",
   775 => x"2e8a3875",
   776 => x"80f82e09",
   777 => x"81068938",
   778 => x"76841871",
   779 => x"085e5854",
   780 => x"7580e42e",
   781 => x"9f387580",
   782 => x"e4268a38",
   783 => x"7580e32e",
   784 => x"be38998a",
   785 => x"047580f3",
   786 => x"2ea33875",
   787 => x"80f82e89",
   788 => x"38998a04",
   789 => x"8a5398db",
   790 => x"049053b4",
   791 => x"a0527b51",
   792 => x"97832db3",
   793 => x"c008b4a0",
   794 => x"5a55999a",
   795 => x"04768418",
   796 => x"71087054",
   797 => x"5b585495",
   798 => x"da2d8055",
   799 => x"999a0476",
   800 => x"84187108",
   801 => x"58585499",
   802 => x"c504a551",
   803 => x"95b82d75",
   804 => x"5195b82d",
   805 => x"82185899",
   806 => x"cd0474ff",
   807 => x"16565480",
   808 => x"7425aa38",
   809 => x"78708105",
   810 => x"5a80f52d",
   811 => x"70525695",
   812 => x"b82d8118",
   813 => x"58999a04",
   814 => x"75a52e09",
   815 => x"81068638",
   816 => x"815e99cd",
   817 => x"04755195",
   818 => x"b82d8118",
   819 => x"58811b5b",
   820 => x"837b25fe",
   821 => x"ac3875fe",
   822 => x"9f387eb3",
   823 => x"c00c0280",
   824 => x"c0050d04",
   825 => x"02ec050d",
   826 => x"76557480",
   827 => x"f52d5170",
   828 => x"802e81f2",
   829 => x"38b4e408",
   830 => x"70828080",
   831 => x"29a9bc08",
   832 => x"05b4e008",
   833 => x"11515252",
   834 => x"718f24de",
   835 => x"38747081",
   836 => x"055680f5",
   837 => x"2d527180",
   838 => x"2e81cb38",
   839 => x"71882e09",
   840 => x"81069c38",
   841 => x"800bb4e0",
   842 => x"0825b838",
   843 => x"ff1151a0",
   844 => x"7181b72d",
   845 => x"b4e008ff",
   846 => x"05b4e00c",
   847 => x"9b8b0471",
   848 => x"8a2e0981",
   849 => x"069d38b4",
   850 => x"e4088105",
   851 => x"b4e40c80",
   852 => x"0bb4e00c",
   853 => x"b4e40882",
   854 => x"808029a9",
   855 => x"bc080551",
   856 => x"9b8b0471",
   857 => x"71708105",
   858 => x"5381b72d",
   859 => x"b4e00881",
   860 => x"05b4e00c",
   861 => x"b4e008a0",
   862 => x"2e098106",
   863 => x"8e38800b",
   864 => x"b4e00cb4",
   865 => x"e4088105",
   866 => x"b4e40c8f",
   867 => x"0bb4e408",
   868 => x"2580c738",
   869 => x"a9bc0882",
   870 => x"80801171",
   871 => x"53555381",
   872 => x"ff527370",
   873 => x"84055508",
   874 => x"71708405",
   875 => x"530cff12",
   876 => x"52718025",
   877 => x"ed388880",
   878 => x"13518f52",
   879 => x"80717084",
   880 => x"05530cff",
   881 => x"12527180",
   882 => x"25f23880",
   883 => x"0bb4e00c",
   884 => x"8f0bb4e4",
   885 => x"0c9e8080",
   886 => x"13518f0b",
   887 => x"b4e40825",
   888 => x"feab3899",
   889 => x"ea040294",
   890 => x"050d0402",
   891 => x"f4050d02",
   892 => x"930580f5",
   893 => x"2d028c05",
   894 => x"81b72d80",
   895 => x"02840589",
   896 => x"0581b72d",
   897 => x"028c05fc",
   898 => x"055199e4",
   899 => x"2d810bb3",
   900 => x"c00c028c",
   901 => x"050d0402",
   902 => x"fc050d72",
   903 => x"5199e42d",
   904 => x"800bb3c0",
   905 => x"0c028405",
   906 => x"0d0402f8",
   907 => x"050da9bc",
   908 => x"08528ffc",
   909 => x"51807270",
   910 => x"8405540c",
   911 => x"fc115170",
   912 => x"8025f238",
   913 => x"0288050d",
   914 => x"0402fc05",
   915 => x"0d725180",
   916 => x"710c800b",
   917 => x"84120c80",
   918 => x"0b88120c",
   919 => x"800b8c12",
   920 => x"0c028405",
   921 => x"0d0402f0",
   922 => x"050d7570",
   923 => x"08841208",
   924 => x"535353ff",
   925 => x"5471712e",
   926 => x"9b388413",
   927 => x"08708429",
   928 => x"14931180",
   929 => x"f52d8416",
   930 => x"08811187",
   931 => x"0684180c",
   932 => x"52565151",
   933 => x"73b3c00c",
   934 => x"0290050d",
   935 => x"0402f405",
   936 => x"0d747008",
   937 => x"84120853",
   938 => x"53537072",
   939 => x"248f3872",
   940 => x"08841408",
   941 => x"71713152",
   942 => x"52529dca",
   943 => x"04720884",
   944 => x"14087171",
   945 => x"31880552",
   946 => x"525271b3",
   947 => x"c00c028c",
   948 => x"050d0402",
   949 => x"f8050da2",
   950 => x"b72da2aa",
   951 => x"2de00870",
   952 => x"8b2a7081",
   953 => x"06515252",
   954 => x"70802e9d",
   955 => x"38b9c808",
   956 => x"708429b9",
   957 => x"d8057381",
   958 => x"ff06710c",
   959 => x"5151b9c8",
   960 => x"08811187",
   961 => x"06b9c80c",
   962 => x"51718a2a",
   963 => x"70810651",
   964 => x"5170802e",
   965 => x"a838b9d0",
   966 => x"08b9d408",
   967 => x"52527171",
   968 => x"2e9b38b9",
   969 => x"d0087084",
   970 => x"29b9f805",
   971 => x"7008e00c",
   972 => x"5151b9d0",
   973 => x"08811187",
   974 => x"06b9d00c",
   975 => x"51a2b12d",
   976 => x"0288050d",
   977 => x"0402f405",
   978 => x"0d74538c",
   979 => x"13088111",
   980 => x"87068815",
   981 => x"08545151",
   982 => x"71712eef",
   983 => x"38a2b72d",
   984 => x"8c130870",
   985 => x"84291477",
   986 => x"b0120c51",
   987 => x"518c1308",
   988 => x"81118706",
   989 => x"8c150c51",
   990 => x"9dd32da2",
   991 => x"b12d028c",
   992 => x"050d0402",
   993 => x"fc050db9",
   994 => x"c8519cc9",
   995 => x"2d9dd351",
   996 => x"a2a62da1",
   997 => x"de2d0284",
   998 => x"050d0402",
   999 => x"e4050d80",
  1000 => x"57a1a904",
  1001 => x"b3c00881",
  1002 => x"f02e0981",
  1003 => x"06893881",
  1004 => x"0bb4f00c",
  1005 => x"a1a904b3",
  1006 => x"c00881e0",
  1007 => x"2e098106",
  1008 => x"8938810b",
  1009 => x"b4f40ca1",
  1010 => x"a904b3c0",
  1011 => x"0854b4f4",
  1012 => x"08802e88",
  1013 => x"38b3c008",
  1014 => x"81800554",
  1015 => x"b4f00881",
  1016 => x"9c38830b",
  1017 => x"a9c01581",
  1018 => x"b72d7480",
  1019 => x"ff24b138",
  1020 => x"b4ec0882",
  1021 => x"2a708106",
  1022 => x"b4e80870",
  1023 => x"872b8180",
  1024 => x"07781182",
  1025 => x"2b515658",
  1026 => x"5154738b",
  1027 => x"38758180",
  1028 => x"29157082",
  1029 => x"2b5153ab",
  1030 => x"c0130853",
  1031 => x"7281b638",
  1032 => x"800bb4f4",
  1033 => x"0c7480d9",
  1034 => x"2e80c738",
  1035 => x"7480d924",
  1036 => x"8f387492",
  1037 => x"2ebc3874",
  1038 => x"80d82e93",
  1039 => x"38a1a404",
  1040 => x"7480f72e",
  1041 => x"a0387480",
  1042 => x"fe2e8f38",
  1043 => x"a1a404b4",
  1044 => x"ec088432",
  1045 => x"b4ec0ca0",
  1046 => x"ed04b4ec",
  1047 => x"088132b4",
  1048 => x"ec0ca0ed",
  1049 => x"04b4ec08",
  1050 => x"8232b4ec",
  1051 => x"0c8157a1",
  1052 => x"a404b4e8",
  1053 => x"088107b4",
  1054 => x"e80ca1a4",
  1055 => x"04a9c014",
  1056 => x"80f52d81",
  1057 => x"fe065372",
  1058 => x"a9c01581",
  1059 => x"b72d7492",
  1060 => x"2e8a3874",
  1061 => x"80d92e09",
  1062 => x"81068938",
  1063 => x"b4e808fe",
  1064 => x"06b4e80c",
  1065 => x"800bb4f0",
  1066 => x"0cb9c851",
  1067 => x"9ce62db3",
  1068 => x"c00855b3",
  1069 => x"c008ff24",
  1070 => x"fdea3876",
  1071 => x"802e9438",
  1072 => x"81ed52b9",
  1073 => x"c8519ec5",
  1074 => x"2db4ec08",
  1075 => x"52b9c851",
  1076 => x"9ec52d80",
  1077 => x"5372b3c0",
  1078 => x"0c029c05",
  1079 => x"0d0402fc",
  1080 => x"050d8051",
  1081 => x"800ba9c0",
  1082 => x"1281b72d",
  1083 => x"81115181",
  1084 => x"ff7125f0",
  1085 => x"38028405",
  1086 => x"0d0402f4",
  1087 => x"050d7451",
  1088 => x"a2b72da9",
  1089 => x"c01180f5",
  1090 => x"2d7081ff",
  1091 => x"0671fd06",
  1092 => x"52545271",
  1093 => x"a9c01281",
  1094 => x"b72da2b1",
  1095 => x"2d72b3c0",
  1096 => x"0c028c05",
  1097 => x"0d047198",
  1098 => x"0c04ffb0",
  1099 => x"08b3c00c",
  1100 => x"04810bff",
  1101 => x"b00c0480",
  1102 => x"0bffb00c",
  1103 => x"0402e805",
  1104 => x"0d787871",
  1105 => x"54575372",
  1106 => x"80258438",
  1107 => x"83135271",
  1108 => x"822cff05",
  1109 => x"5372ff2e",
  1110 => x"80c03875",
  1111 => x"70840557",
  1112 => x"08548755",
  1113 => x"739c2ab0",
  1114 => x"0552b972",
  1115 => x"27843887",
  1116 => x"12527151",
  1117 => x"95b82d73",
  1118 => x"842bff16",
  1119 => x"56547480",
  1120 => x"25e238a0",
  1121 => x"5195b82d",
  1122 => x"72870652",
  1123 => x"7186388a",
  1124 => x"5195b82d",
  1125 => x"ff1353a2",
  1126 => x"d5048a51",
  1127 => x"95b82d02",
  1128 => x"98050d04",
  1129 => x"b3cc0802",
  1130 => x"b3cc0cff",
  1131 => x"3d0d800b",
  1132 => x"b3cc08fc",
  1133 => x"050cb3cc",
  1134 => x"08880508",
  1135 => x"8106ff11",
  1136 => x"700970b3",
  1137 => x"cc088c05",
  1138 => x"0806b3cc",
  1139 => x"08fc0508",
  1140 => x"11b3cc08",
  1141 => x"fc050cb3",
  1142 => x"cc088805",
  1143 => x"08812ab3",
  1144 => x"cc088805",
  1145 => x"0cb3cc08",
  1146 => x"8c050810",
  1147 => x"b3cc088c",
  1148 => x"050c5151",
  1149 => x"5151b3cc",
  1150 => x"08880508",
  1151 => x"802e8438",
  1152 => x"ffb439b3",
  1153 => x"cc08fc05",
  1154 => x"0870b3c0",
  1155 => x"0c51833d",
  1156 => x"0db3cc0c",
  1157 => x"04000000",
  1158 => x"00ffffff",
  1159 => x"ff00ffff",
  1160 => x"ffff00ff",
  1161 => x"ffffff00",
  1162 => x"496e6974",
  1163 => x"69616c69",
  1164 => x"7a696e67",
  1165 => x"20534420",
  1166 => x"63617264",
  1167 => x"0a000000",
  1168 => x"4d535833",
  1169 => x"42494f53",
  1170 => x"53595300",
  1171 => x"42494f53",
  1172 => x"5f4d3250",
  1173 => x"524f4d00",
  1174 => x"4f70656e",
  1175 => x"65642066",
  1176 => x"696c652c",
  1177 => x"206c6f61",
  1178 => x"64696e67",
  1179 => x"2e2e2e0a",
  1180 => x"00000000",
  1181 => x"52656164",
  1182 => x"20626c6f",
  1183 => x"636b2066",
  1184 => x"61696c65",
  1185 => x"640a0000",
  1186 => x"4c6f6164",
  1187 => x"696e6720",
  1188 => x"42494f53",
  1189 => x"20666169",
  1190 => x"6c65640a",
  1191 => x"00000000",
  1192 => x"52656164",
  1193 => x"696e6720",
  1194 => x"4d42520a",
  1195 => x"00000000",
  1196 => x"52656164",
  1197 => x"206f6620",
  1198 => x"4d425220",
  1199 => x"6661696c",
  1200 => x"65640a00",
  1201 => x"4d425220",
  1202 => x"73756363",
  1203 => x"65737366",
  1204 => x"756c6c79",
  1205 => x"20726561",
  1206 => x"640a0000",
  1207 => x"46415431",
  1208 => x"36202020",
  1209 => x"00000000",
  1210 => x"46415433",
  1211 => x"32202020",
  1212 => x"00000000",
  1213 => x"50617274",
  1214 => x"6974696f",
  1215 => x"6e636f75",
  1216 => x"6e742025",
  1217 => x"640a0000",
  1218 => x"4e6f2070",
  1219 => x"61727469",
  1220 => x"74696f6e",
  1221 => x"20736967",
  1222 => x"6e617475",
  1223 => x"72652066",
  1224 => x"6f756e64",
  1225 => x"0a000000",
  1226 => x"52656164",
  1227 => x"696e6720",
  1228 => x"626f6f74",
  1229 => x"20736563",
  1230 => x"746f7220",
  1231 => x"25640a00",
  1232 => x"52656164",
  1233 => x"20626f6f",
  1234 => x"74207365",
  1235 => x"63746f72",
  1236 => x"2066726f",
  1237 => x"6d206669",
  1238 => x"72737420",
  1239 => x"70617274",
  1240 => x"6974696f",
  1241 => x"6e0a0000",
  1242 => x"48756e74",
  1243 => x"696e6720",
  1244 => x"666f7220",
  1245 => x"66696c65",
  1246 => x"73797374",
  1247 => x"656d0a00",
  1248 => x"556e7375",
  1249 => x"70706f72",
  1250 => x"74656420",
  1251 => x"70617274",
  1252 => x"6974696f",
  1253 => x"6e207479",
  1254 => x"7065210d",
  1255 => x"00000000",
  1256 => x"436c7573",
  1257 => x"74657220",
  1258 => x"73697a65",
  1259 => x"3a202564",
  1260 => x"2c20436c",
  1261 => x"75737465",
  1262 => x"72206d61",
  1263 => x"736b2c20",
  1264 => x"25640a00",
  1265 => x"47657443",
  1266 => x"6c757374",
  1267 => x"65722072",
  1268 => x"65616469",
  1269 => x"6e672073",
  1270 => x"6563746f",
  1271 => x"72202564",
  1272 => x"0a000000",
  1273 => x"52656164",
  1274 => x"696e6720",
  1275 => x"64697265",
  1276 => x"63746f72",
  1277 => x"79207365",
  1278 => x"63746f72",
  1279 => x"2025640a",
  1280 => x"00000000",
  1281 => x"47657446",
  1282 => x"41544c69",
  1283 => x"6e6b2072",
  1284 => x"65747572",
  1285 => x"6e656420",
  1286 => x"25640a00",
  1287 => x"436d645f",
  1288 => x"696e6974",
  1289 => x"0a000000",
  1290 => x"636d645f",
  1291 => x"434d4438",
  1292 => x"20726573",
  1293 => x"706f6e73",
  1294 => x"653a2025",
  1295 => x"640a0000",
  1296 => x"434d4438",
  1297 => x"5f342072",
  1298 => x"6573706f",
  1299 => x"6e73653a",
  1300 => x"2025640a",
  1301 => x"00000000",
  1302 => x"53444843",
  1303 => x"20496e69",
  1304 => x"7469616c",
  1305 => x"697a6174",
  1306 => x"696f6e20",
  1307 => x"6572726f",
  1308 => x"72210a00",
  1309 => x"434d4435",
  1310 => x"38202564",
  1311 => x"0a202000",
  1312 => x"434d4435",
  1313 => x"385f3220",
  1314 => x"25640a20",
  1315 => x"20000000",
  1316 => x"53504920",
  1317 => x"496e6974",
  1318 => x"28290a00",
  1319 => x"52656164",
  1320 => x"20636f6d",
  1321 => x"6d616e64",
  1322 => x"20666169",
  1323 => x"6c656420",
  1324 => x"61742025",
  1325 => x"64202825",
  1326 => x"64290a00",
  1327 => x"ffffe000",
  1328 => x"00000000",
  1329 => x"00000000",
  1330 => x"00000000",
  1331 => x"00000000",
  1332 => x"00000000",
  1333 => x"00000000",
  1334 => x"00000000",
  1335 => x"00000000",
  1336 => x"00000000",
  1337 => x"00000000",
  1338 => x"00000000",
  1339 => x"00000000",
  1340 => x"00000000",
  1341 => x"00000000",
  1342 => x"00000000",
  1343 => x"00000000",
  1344 => x"00000000",
  1345 => x"00000000",
  1346 => x"00000000",
  1347 => x"00000000",
  1348 => x"00000000",
  1349 => x"00000000",
  1350 => x"00000000",
  1351 => x"00000000",
  1352 => x"00000000",
  1353 => x"00000000",
  1354 => x"00000000",
  1355 => x"00000000",
  1356 => x"00000000",
  1357 => x"00000000",
  1358 => x"00000000",
  1359 => x"00000000",
  1360 => x"00000000",
  1361 => x"00000000",
  1362 => x"00000000",
  1363 => x"00000000",
  1364 => x"00000000",
  1365 => x"00000000",
  1366 => x"00000000",
  1367 => x"00000000",
  1368 => x"00000000",
  1369 => x"00000000",
  1370 => x"00000000",
  1371 => x"00000000",
  1372 => x"00000000",
  1373 => x"00000000",
  1374 => x"00000000",
  1375 => x"00000000",
  1376 => x"00000000",
  1377 => x"00000000",
  1378 => x"00000000",
  1379 => x"00000000",
  1380 => x"00000000",
  1381 => x"00000000",
  1382 => x"00000000",
  1383 => x"00000000",
  1384 => x"00000000",
  1385 => x"00000000",
  1386 => x"00000000",
  1387 => x"00000000",
  1388 => x"00000000",
  1389 => x"00000000",
  1390 => x"00000000",
  1391 => x"00000000",
  1392 => x"00000000",
  1393 => x"00000000",
  1394 => x"00000000",
  1395 => x"00000000",
  1396 => x"00000000",
  1397 => x"00000000",
  1398 => x"00000000",
  1399 => x"00000000",
  1400 => x"00000000",
  1401 => x"00000000",
  1402 => x"00000000",
  1403 => x"00000000",
  1404 => x"00000000",
  1405 => x"00000009",
  1406 => x"00000000",
  1407 => x"00000000",
  1408 => x"00000000",
  1409 => x"00000000",
  1410 => x"00000000",
  1411 => x"00000000",
  1412 => x"00000000",
  1413 => x"00000071",
  1414 => x"00000031",
  1415 => x"00000000",
  1416 => x"00000000",
  1417 => x"00000000",
  1418 => x"0000007a",
  1419 => x"00000073",
  1420 => x"00000061",
  1421 => x"00000077",
  1422 => x"00000032",
  1423 => x"00000000",
  1424 => x"00000000",
  1425 => x"00000063",
  1426 => x"00000078",
  1427 => x"00000064",
  1428 => x"00000065",
  1429 => x"00000034",
  1430 => x"00000033",
  1431 => x"00000000",
  1432 => x"00000000",
  1433 => x"00000020",
  1434 => x"00000076",
  1435 => x"00000066",
  1436 => x"00000074",
  1437 => x"00000072",
  1438 => x"00000035",
  1439 => x"00000000",
  1440 => x"00000000",
  1441 => x"0000006e",
  1442 => x"00000062",
  1443 => x"00000068",
  1444 => x"00000067",
  1445 => x"00000079",
  1446 => x"00000036",
  1447 => x"00000000",
  1448 => x"00000000",
  1449 => x"00000000",
  1450 => x"0000006d",
  1451 => x"0000006a",
  1452 => x"00000075",
  1453 => x"00000037",
  1454 => x"00000038",
  1455 => x"00000000",
  1456 => x"00000000",
  1457 => x"0000002c",
  1458 => x"0000006b",
  1459 => x"00000069",
  1460 => x"0000006f",
  1461 => x"00000030",
  1462 => x"00000039",
  1463 => x"00000000",
  1464 => x"00000000",
  1465 => x"0000002e",
  1466 => x"0000002f",
  1467 => x"0000006c",
  1468 => x"0000003b",
  1469 => x"00000070",
  1470 => x"0000002d",
  1471 => x"00000000",
  1472 => x"00000000",
  1473 => x"00000000",
  1474 => x"00000027",
  1475 => x"00000000",
  1476 => x"0000005b",
  1477 => x"0000003d",
  1478 => x"00000000",
  1479 => x"00000000",
  1480 => x"00000000",
  1481 => x"00000000",
  1482 => x"0000000a",
  1483 => x"0000005d",
  1484 => x"00000000",
  1485 => x"00000023",
  1486 => x"00000000",
  1487 => x"00000000",
  1488 => x"00000000",
  1489 => x"00000000",
  1490 => x"00000000",
  1491 => x"00000000",
  1492 => x"00000000",
  1493 => x"00000000",
  1494 => x"00000008",
  1495 => x"00000000",
  1496 => x"00000000",
  1497 => x"00000031",
  1498 => x"00000000",
  1499 => x"00000034",
  1500 => x"00000037",
  1501 => x"00000000",
  1502 => x"00000000",
  1503 => x"00000000",
  1504 => x"00000030",
  1505 => x"0000002e",
  1506 => x"00000032",
  1507 => x"00000035",
  1508 => x"00000036",
  1509 => x"00000038",
  1510 => x"0000001b",
  1511 => x"00000000",
  1512 => x"00000000",
  1513 => x"0000002b",
  1514 => x"00000033",
  1515 => x"00000000",
  1516 => x"0000002a",
  1517 => x"00000039",
  1518 => x"00000000",
  1519 => x"00000000",
  1520 => x"00000000",
  1521 => x"00000000",
  1522 => x"00000000",
  1523 => x"00000000",
  1524 => x"00000000",
  1525 => x"00000000",
  1526 => x"00000000",
  1527 => x"00000000",
  1528 => x"00000000",
  1529 => x"00000000",
  1530 => x"00000000",
  1531 => x"00000000",
  1532 => x"00000000",
  1533 => x"00000008",
  1534 => x"00000000",
  1535 => x"00000000",
  1536 => x"00000000",
  1537 => x"00000000",
  1538 => x"00000000",
  1539 => x"00000000",
  1540 => x"00000000",
  1541 => x"00000051",
  1542 => x"00000021",
  1543 => x"00000000",
  1544 => x"00000000",
  1545 => x"00000000",
  1546 => x"0000005a",
  1547 => x"00000053",
  1548 => x"00000041",
  1549 => x"00000057",
  1550 => x"00000022",
  1551 => x"00000000",
  1552 => x"00000000",
  1553 => x"00000043",
  1554 => x"00000058",
  1555 => x"00000044",
  1556 => x"00000045",
  1557 => x"00000024",
  1558 => x"000000a3",
  1559 => x"00000000",
  1560 => x"00000000",
  1561 => x"00000020",
  1562 => x"00000056",
  1563 => x"00000046",
  1564 => x"00000054",
  1565 => x"00000052",
  1566 => x"00000025",
  1567 => x"00000000",
  1568 => x"00000000",
  1569 => x"0000004e",
  1570 => x"00000042",
  1571 => x"00000048",
  1572 => x"00000047",
  1573 => x"00000059",
  1574 => x"0000005e",
  1575 => x"00000000",
  1576 => x"00000000",
  1577 => x"00000000",
  1578 => x"0000004d",
  1579 => x"0000004a",
  1580 => x"00000055",
  1581 => x"00000026",
  1582 => x"0000002a",
  1583 => x"00000000",
  1584 => x"00000000",
  1585 => x"0000003c",
  1586 => x"0000004b",
  1587 => x"00000049",
  1588 => x"0000004f",
  1589 => x"00000029",
  1590 => x"00000028",
  1591 => x"00000000",
  1592 => x"00000000",
  1593 => x"0000003e",
  1594 => x"0000003f",
  1595 => x"0000004c",
  1596 => x"0000003a",
  1597 => x"00000050",
  1598 => x"0000005f",
  1599 => x"00000000",
  1600 => x"00000000",
  1601 => x"00000000",
  1602 => x"0000003f",
  1603 => x"00000000",
  1604 => x"0000007b",
  1605 => x"0000002b",
  1606 => x"00000000",
  1607 => x"00000000",
  1608 => x"00000000",
  1609 => x"00000000",
  1610 => x"0000000a",
  1611 => x"0000007d",
  1612 => x"00000000",
  1613 => x"0000007e",
  1614 => x"00000000",
  1615 => x"00000000",
  1616 => x"00000000",
  1617 => x"00000000",
  1618 => x"00000000",
  1619 => x"00000000",
  1620 => x"00000000",
  1621 => x"00000000",
  1622 => x"00000009",
  1623 => x"00000000",
  1624 => x"00000000",
  1625 => x"00000031",
  1626 => x"00000000",
  1627 => x"00000034",
  1628 => x"00000037",
  1629 => x"00000000",
  1630 => x"00000000",
  1631 => x"00000000",
  1632 => x"00000030",
  1633 => x"0000002e",
  1634 => x"00000032",
  1635 => x"00000035",
  1636 => x"00000036",
  1637 => x"00000038",
  1638 => x"0000001b",
  1639 => x"00000000",
  1640 => x"00000000",
  1641 => x"0000002b",
  1642 => x"00000033",
  1643 => x"00000000",
  1644 => x"0000002a",
  1645 => x"00000039",
  1646 => x"00000000",
  1647 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

