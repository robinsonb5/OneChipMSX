-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b0bb3",
     9 => x"e0080b0b",
    10 => x"0bb3e408",
    11 => x"0b0b0bb3",
    12 => x"e8080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"b3e80c0b",
    16 => x"0b0bb3e4",
    17 => x"0c0b0b0b",
    18 => x"b3e00c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0ba48c",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"b3e070ba",
    57 => x"b8278b38",
    58 => x"80717084",
    59 => x"05530c81",
    60 => x"e2048c51",
    61 => x"81f70402",
    62 => x"d8050d81",
    63 => x"0bfec40c",
    64 => x"b90bfec0",
    65 => x"0c840bfe",
    66 => x"c40ca49c",
    67 => x"5195ce2d",
    68 => x"9ef72da2",
    69 => x"a52da4bc",
    70 => x"5195ce2d",
    71 => x"92ef2db3",
    72 => x"e008802e",
    73 => x"81c538a4",
    74 => x"d45195ce",
    75 => x"2d84c22d",
    76 => x"a4ec52b5",
    77 => x"98518b97",
    78 => x"2db3e008",
    79 => x"81ff0653",
    80 => x"72802e81",
    81 => x"a038a4f8",
    82 => x"5195ce2d",
    83 => x"b59c0857",
    84 => x"80597877",
    85 => x"25819438",
    86 => x"b5b052b5",
    87 => x"98518dee",
    88 => x"2db3e008",
    89 => x"81ff06b5",
    90 => x"b05b5380",
    91 => x"5872782e",
    92 => x"098106b1",
    93 => x"3883b804",
    94 => x"79708405",
    95 => x"5b087081",
    96 => x"ff067188",
    97 => x"2c7081ff",
    98 => x"0673902c",
    99 => x"7081ff06",
   100 => x"75982afe",
   101 => x"c80cfec8",
   102 => x"0c58fec8",
   103 => x"0c57fec8",
   104 => x"0c841959",
   105 => x"53765384",
   106 => x"80772584",
   107 => x"38848053",
   108 => x"727824c4",
   109 => x"3883be04",
   110 => x"a5945195",
   111 => x"ce2db598",
   112 => x"518dc12d",
   113 => x"fc801781",
   114 => x"1a5a57ae",
   115 => x"5195ac2d",
   116 => x"78bf0653",
   117 => x"7286388a",
   118 => x"5195ac2d",
   119 => x"768024fe",
   120 => x"f73883eb",
   121 => x"04a5a851",
   122 => x"95ce2d82",
   123 => x"0bfec40c",
   124 => x"9f8f2db3",
   125 => x"e008802e",
   126 => x"f738b3e0",
   127 => x"085195ac",
   128 => x"2d83f004",
   129 => x"02e8050d",
   130 => x"77797b58",
   131 => x"55558053",
   132 => x"727625a3",
   133 => x"38747081",
   134 => x"055680f5",
   135 => x"2d747081",
   136 => x"055680f5",
   137 => x"2d525271",
   138 => x"712e8638",
   139 => x"815184b9",
   140 => x"04811353",
   141 => x"84900480",
   142 => x"5170b3e0",
   143 => x"0c029805",
   144 => x"0d0402d8",
   145 => x"050d800b",
   146 => x"b9c80ca5",
   147 => x"c05195ce",
   148 => x"2db5b052",
   149 => x"80519489",
   150 => x"2db3e008",
   151 => x"54b3e008",
   152 => x"8c38a5d0",
   153 => x"5195ce2d",
   154 => x"73558a95",
   155 => x"04a5e451",
   156 => x"95ce2d80",
   157 => x"56810bb5",
   158 => x"a40c8853",
   159 => x"a5fc52b5",
   160 => x"e6518484",
   161 => x"2db3e008",
   162 => x"762e0981",
   163 => x"068738b3",
   164 => x"e008b5a4",
   165 => x"0c8853a6",
   166 => x"8852b682",
   167 => x"5184842d",
   168 => x"b3e00887",
   169 => x"38b3e008",
   170 => x"b5a40cb5",
   171 => x"a40852a6",
   172 => x"945197d6",
   173 => x"2db5a408",
   174 => x"802e8187",
   175 => x"38b8f60b",
   176 => x"80f52db8",
   177 => x"f70b80f5",
   178 => x"2d71982b",
   179 => x"71902b07",
   180 => x"b8f80b80",
   181 => x"f52d7088",
   182 => x"2b7207b8",
   183 => x"f90b80f5",
   184 => x"2d7107b9",
   185 => x"ae0b80f5",
   186 => x"2db9af0b",
   187 => x"80f52d71",
   188 => x"882b0753",
   189 => x"5f54525a",
   190 => x"56575573",
   191 => x"81abaa2e",
   192 => x"0981068d",
   193 => x"38755196",
   194 => x"962db3e0",
   195 => x"085686a1",
   196 => x"047382d4",
   197 => x"d52e8a38",
   198 => x"a6a85195",
   199 => x"ce2d87d6",
   200 => x"047552a6",
   201 => x"c85197d6",
   202 => x"2db5b052",
   203 => x"75519489",
   204 => x"2db3e008",
   205 => x"55b3e008",
   206 => x"802e83d9",
   207 => x"38a6e051",
   208 => x"95ce2da7",
   209 => x"885197d6",
   210 => x"2d8853a6",
   211 => x"8852b682",
   212 => x"5184842d",
   213 => x"b3e00889",
   214 => x"38810bb9",
   215 => x"c80c86fc",
   216 => x"048853a5",
   217 => x"fc52b5e6",
   218 => x"5184842d",
   219 => x"b3e00880",
   220 => x"2e8a38a7",
   221 => x"a05197d6",
   222 => x"2d87d604",
   223 => x"b9ae0b80",
   224 => x"f52d5473",
   225 => x"80d52e09",
   226 => x"810680ca",
   227 => x"38b9af0b",
   228 => x"80f52d54",
   229 => x"7381aa2e",
   230 => x"098106ba",
   231 => x"38800bb5",
   232 => x"b00b80f5",
   233 => x"2d565474",
   234 => x"81e92e83",
   235 => x"38815474",
   236 => x"81eb2e8c",
   237 => x"38805573",
   238 => x"752e0981",
   239 => x"0682d638",
   240 => x"b5bb0b80",
   241 => x"f52d5978",
   242 => x"8d38b5bc",
   243 => x"0b80f52d",
   244 => x"5473822e",
   245 => x"86388055",
   246 => x"8a9504b5",
   247 => x"bd0b80f5",
   248 => x"2d70b9d0",
   249 => x"0cff1170",
   250 => x"b9c40c54",
   251 => x"52a7c051",
   252 => x"97d62db5",
   253 => x"be0b80f5",
   254 => x"2db5bf0b",
   255 => x"80f52d56",
   256 => x"76057582",
   257 => x"80290570",
   258 => x"b9b80cb5",
   259 => x"c00b80f5",
   260 => x"2d70b9b4",
   261 => x"0cb9c808",
   262 => x"59575876",
   263 => x"802e81a5",
   264 => x"388853a6",
   265 => x"8852b682",
   266 => x"5184842d",
   267 => x"7855b3e0",
   268 => x"0881e238",
   269 => x"b9d00870",
   270 => x"842bb9b0",
   271 => x"0c70b9cc",
   272 => x"0cb5d50b",
   273 => x"80f52db5",
   274 => x"d40b80f5",
   275 => x"2d718280",
   276 => x"2905b5d6",
   277 => x"0b80f52d",
   278 => x"70848080",
   279 => x"2912b5d7",
   280 => x"0b80f52d",
   281 => x"7081800a",
   282 => x"291270b5",
   283 => x"a80cb9b4",
   284 => x"087129b9",
   285 => x"b8080570",
   286 => x"b9d80cb5",
   287 => x"dd0b80f5",
   288 => x"2db5dc0b",
   289 => x"80f52d71",
   290 => x"82802905",
   291 => x"b5de0b80",
   292 => x"f52d7084",
   293 => x"80802912",
   294 => x"b5df0b80",
   295 => x"f52d7098",
   296 => x"2b81f00a",
   297 => x"06720570",
   298 => x"b5ac0cfe",
   299 => x"117e2977",
   300 => x"05b9c00c",
   301 => x"52575257",
   302 => x"5d575152",
   303 => x"5f525c57",
   304 => x"57578a93",
   305 => x"04b5c20b",
   306 => x"80f52db5",
   307 => x"c10b80f5",
   308 => x"2d718280",
   309 => x"290570b9",
   310 => x"b00c70a0",
   311 => x"2983ff05",
   312 => x"70892a70",
   313 => x"b9cc0cb5",
   314 => x"c70b80f5",
   315 => x"2db5c60b",
   316 => x"80f52d71",
   317 => x"82802905",
   318 => x"70b5a80c",
   319 => x"7b71291e",
   320 => x"70b9c00c",
   321 => x"7db5ac0c",
   322 => x"7305b9d8",
   323 => x"0c555e51",
   324 => x"51555581",
   325 => x"5574b3e0",
   326 => x"0c02a805",
   327 => x"0d0402ec",
   328 => x"050d7670",
   329 => x"872c7180",
   330 => x"ff065755",
   331 => x"53b9c808",
   332 => x"8a387288",
   333 => x"2c7381ff",
   334 => x"065654b9",
   335 => x"b8081452",
   336 => x"a7e45197",
   337 => x"d62db5b0",
   338 => x"52b9b808",
   339 => x"14519489",
   340 => x"2db3e008",
   341 => x"53b3e008",
   342 => x"802eb338",
   343 => x"b9c80880",
   344 => x"2e983874",
   345 => x"8429b5b0",
   346 => x"05700852",
   347 => x"5396962d",
   348 => x"b3e008f0",
   349 => x"0a06558b",
   350 => x"8c047410",
   351 => x"b5b00570",
   352 => x"80e02d52",
   353 => x"5396c62d",
   354 => x"b3e00855",
   355 => x"745372b3",
   356 => x"e00c0294",
   357 => x"050d0402",
   358 => x"c8050d7f",
   359 => x"615f5c80",
   360 => x"0bb5ac08",
   361 => x"b9c00859",
   362 => x"5956b9c8",
   363 => x"08762e8a",
   364 => x"38b9d008",
   365 => x"842b598b",
   366 => x"c004b9cc",
   367 => x"08842b59",
   368 => x"805a7979",
   369 => x"2781b638",
   370 => x"798f06a0",
   371 => x"17575473",
   372 => x"97387652",
   373 => x"a8845197",
   374 => x"d62db5b0",
   375 => x"52765181",
   376 => x"17579489",
   377 => x"2db5b056",
   378 => x"807680f5",
   379 => x"2d565474",
   380 => x"742e8338",
   381 => x"81547481",
   382 => x"e52e80fb",
   383 => x"38817075",
   384 => x"06555d73",
   385 => x"802e80ef",
   386 => x"388b1680",
   387 => x"f52d9806",
   388 => x"5b7a80e3",
   389 => x"38755195",
   390 => x"ce2d8b53",
   391 => x"7d527551",
   392 => x"84842db3",
   393 => x"e00880cf",
   394 => x"389c1608",
   395 => x"5196962d",
   396 => x"b3e00884",
   397 => x"1d0c9a16",
   398 => x"80e02d51",
   399 => x"96c62db3",
   400 => x"e008b3e0",
   401 => x"08881e0c",
   402 => x"b3e00855",
   403 => x"55b9c808",
   404 => x"802e9838",
   405 => x"941680e0",
   406 => x"2d5196c6",
   407 => x"2db3e008",
   408 => x"902b83ff",
   409 => x"f00a0670",
   410 => x"16515473",
   411 => x"881d0c7a",
   412 => x"7c0c7c54",
   413 => x"8db80481",
   414 => x"1a5a8bc2",
   415 => x"04b9c808",
   416 => x"802eb338",
   417 => x"77518a9e",
   418 => x"2db3e008",
   419 => x"b3e00853",
   420 => x"a8a45258",
   421 => x"97d62d77",
   422 => x"80ffffff",
   423 => x"f8065473",
   424 => x"80ffffff",
   425 => x"f82e8f38",
   426 => x"fe18b9d0",
   427 => x"0829b9d8",
   428 => x"0805578b",
   429 => x"c0048054",
   430 => x"73b3e00c",
   431 => x"02b8050d",
   432 => x"0402f405",
   433 => x"0d747008",
   434 => x"8105710c",
   435 => x"7008b9c4",
   436 => x"08065353",
   437 => x"718e3888",
   438 => x"1308518a",
   439 => x"9e2db3e0",
   440 => x"0888140c",
   441 => x"810bb3e0",
   442 => x"0c028c05",
   443 => x"0d0402f0",
   444 => x"050d7588",
   445 => x"1108fe05",
   446 => x"b9d00829",
   447 => x"b9d80811",
   448 => x"7208b9c4",
   449 => x"08060579",
   450 => x"55535454",
   451 => x"94892db3",
   452 => x"e00853b3",
   453 => x"e008802e",
   454 => x"83388153",
   455 => x"72b3e00c",
   456 => x"0290050d",
   457 => x"0402f405",
   458 => x"0dd45281",
   459 => x"ff720c71",
   460 => x"085381ff",
   461 => x"720c7288",
   462 => x"2b83fe80",
   463 => x"06720870",
   464 => x"81ff0651",
   465 => x"525381ff",
   466 => x"720c7271",
   467 => x"07882b72",
   468 => x"087081ff",
   469 => x"06515253",
   470 => x"81ff720c",
   471 => x"72710788",
   472 => x"2b720870",
   473 => x"81ff0672",
   474 => x"07b3e00c",
   475 => x"5253028c",
   476 => x"050d0402",
   477 => x"f4050d74",
   478 => x"767181ff",
   479 => x"06d40c53",
   480 => x"53b9dc08",
   481 => x"85387189",
   482 => x"2b527198",
   483 => x"2ad40c71",
   484 => x"902a7081",
   485 => x"ff06d40c",
   486 => x"5171882a",
   487 => x"7081ff06",
   488 => x"d40c5171",
   489 => x"81ff06d4",
   490 => x"0c72902a",
   491 => x"7081ff06",
   492 => x"d40c51d4",
   493 => x"087081ff",
   494 => x"06515182",
   495 => x"b8bf5270",
   496 => x"81ff2e09",
   497 => x"81069438",
   498 => x"81ff0bd4",
   499 => x"0cd40870",
   500 => x"81ff06ff",
   501 => x"14545151",
   502 => x"71e53870",
   503 => x"b3e00c02",
   504 => x"8c050d04",
   505 => x"02fc050d",
   506 => x"81c75181",
   507 => x"ff0bd40c",
   508 => x"ff115170",
   509 => x"8025f438",
   510 => x"0284050d",
   511 => x"0402f005",
   512 => x"0d8fe42d",
   513 => x"819c9f53",
   514 => x"805287fc",
   515 => x"80f7518e",
   516 => x"f32db3e0",
   517 => x"0854b3e0",
   518 => x"08812e09",
   519 => x"8106a338",
   520 => x"81ff0bd4",
   521 => x"0c820a52",
   522 => x"849c80e9",
   523 => x"518ef32d",
   524 => x"b3e0088b",
   525 => x"3881ff0b",
   526 => x"d40c7353",
   527 => x"90c8048f",
   528 => x"e42dff13",
   529 => x"5372c138",
   530 => x"72b3e00c",
   531 => x"0290050d",
   532 => x"0402f405",
   533 => x"0d81ff0b",
   534 => x"d40ca8bc",
   535 => x"5195ce2d",
   536 => x"93538052",
   537 => x"87fc80c1",
   538 => x"518ef32d",
   539 => x"b3e0088b",
   540 => x"3881ff0b",
   541 => x"d40c8153",
   542 => x"9184048f",
   543 => x"e42dff13",
   544 => x"5372df38",
   545 => x"72b3e00c",
   546 => x"028c050d",
   547 => x"0402f005",
   548 => x"0d8fe42d",
   549 => x"83aa5284",
   550 => x"9c80c851",
   551 => x"8ef32db3",
   552 => x"e008b3e0",
   553 => x"0853a8c8",
   554 => x"525397d6",
   555 => x"2d72812e",
   556 => x"0981069c",
   557 => x"388ea52d",
   558 => x"b3e00883",
   559 => x"ffff0653",
   560 => x"7283aa2e",
   561 => x"a138b3e0",
   562 => x"0852a8e0",
   563 => x"5197d62d",
   564 => x"90d12d91",
   565 => x"e1048154",
   566 => x"92e604a8",
   567 => x"f85197d6",
   568 => x"2d805492",
   569 => x"e60481ff",
   570 => x"0bd40cb1",
   571 => x"538ffd2d",
   572 => x"b3e00880",
   573 => x"2e80e038",
   574 => x"805287fc",
   575 => x"80fa518e",
   576 => x"f32db3e0",
   577 => x"0880c638",
   578 => x"b3e00852",
   579 => x"a9945197",
   580 => x"d62d81ff",
   581 => x"0bd40cd4",
   582 => x"087081ff",
   583 => x"067054a9",
   584 => x"a0535153",
   585 => x"97d62d81",
   586 => x"ff0bd40c",
   587 => x"81ff0bd4",
   588 => x"0c81ff0b",
   589 => x"d40c81ff",
   590 => x"0bd40c72",
   591 => x"862a7081",
   592 => x"06705651",
   593 => x"5372802e",
   594 => x"9d3891d6",
   595 => x"04b3e008",
   596 => x"52a99451",
   597 => x"97d62d72",
   598 => x"822efeff",
   599 => x"38ff1353",
   600 => x"72ff8a38",
   601 => x"725473b3",
   602 => x"e00c0290",
   603 => x"050d0402",
   604 => x"f4050d81",
   605 => x"0bb9dc0c",
   606 => x"d008708f",
   607 => x"2a708106",
   608 => x"51515372",
   609 => x"f33872d0",
   610 => x"0c8fe42d",
   611 => x"a9b05195",
   612 => x"ce2dd008",
   613 => x"708f2a70",
   614 => x"81065151",
   615 => x"5372f338",
   616 => x"810bd00c",
   617 => x"87538052",
   618 => x"84d480c0",
   619 => x"518ef32d",
   620 => x"b3e00881",
   621 => x"2e943872",
   622 => x"822e0981",
   623 => x"06863880",
   624 => x"5393fa04",
   625 => x"ff135372",
   626 => x"dd38918d",
   627 => x"2db3e008",
   628 => x"b9dc0c81",
   629 => x"5287fc80",
   630 => x"d0518ef3",
   631 => x"2d81ff0b",
   632 => x"d40cd008",
   633 => x"708f2a70",
   634 => x"81065151",
   635 => x"5372f338",
   636 => x"72d00c81",
   637 => x"ff0bd40c",
   638 => x"815372b3",
   639 => x"e00c028c",
   640 => x"050d0480",
   641 => x"0bb3e00c",
   642 => x"0402e005",
   643 => x"0d797b57",
   644 => x"57805881",
   645 => x"ff0bd40c",
   646 => x"d008708f",
   647 => x"2a708106",
   648 => x"51515473",
   649 => x"f3388281",
   650 => x"0bd00c81",
   651 => x"ff0bd40c",
   652 => x"765287fc",
   653 => x"80d1518e",
   654 => x"f32d80db",
   655 => x"c6df55b3",
   656 => x"e008802e",
   657 => x"9038b3e0",
   658 => x"08537652",
   659 => x"a9bc5197",
   660 => x"d62d95a3",
   661 => x"0481ff0b",
   662 => x"d40cd408",
   663 => x"7081ff06",
   664 => x"51547381",
   665 => x"fe2e0981",
   666 => x"069d3880",
   667 => x"ff548ea5",
   668 => x"2db3e008",
   669 => x"76708405",
   670 => x"580cff14",
   671 => x"54738025",
   672 => x"ed388158",
   673 => x"958d04ff",
   674 => x"155574c9",
   675 => x"3881ff0b",
   676 => x"d40cd008",
   677 => x"708f2a70",
   678 => x"81065151",
   679 => x"5473f338",
   680 => x"73d00c77",
   681 => x"b3e00c02",
   682 => x"a0050d04",
   683 => x"02f8050d",
   684 => x"7352c008",
   685 => x"70882a70",
   686 => x"81065151",
   687 => x"5170802e",
   688 => x"f13871c0",
   689 => x"0c71b3e0",
   690 => x"0c028805",
   691 => x"0d0402e8",
   692 => x"050d8078",
   693 => x"57557570",
   694 => x"84055708",
   695 => x"53805472",
   696 => x"982a7388",
   697 => x"2b545271",
   698 => x"802ea238",
   699 => x"c0087088",
   700 => x"2a708106",
   701 => x"51515170",
   702 => x"802ef138",
   703 => x"71c00c81",
   704 => x"15811555",
   705 => x"55837425",
   706 => x"d63871ca",
   707 => x"3874b3e0",
   708 => x"0c029805",
   709 => x"0d0402f4",
   710 => x"050d7470",
   711 => x"882a83fe",
   712 => x"80067072",
   713 => x"982a0772",
   714 => x"882b87fc",
   715 => x"80800673",
   716 => x"982b81f0",
   717 => x"0a067173",
   718 => x"0707b3e0",
   719 => x"0c565153",
   720 => x"51028c05",
   721 => x"0d0402f8",
   722 => x"050d028e",
   723 => x"0580f52d",
   724 => x"74882b07",
   725 => x"7083ffff",
   726 => x"06b3e00c",
   727 => x"51028805",
   728 => x"0d0402f8",
   729 => x"050d7370",
   730 => x"902b7190",
   731 => x"2a07b3e0",
   732 => x"0c520288",
   733 => x"050d0402",
   734 => x"ec050d76",
   735 => x"53805572",
   736 => x"75258b38",
   737 => x"ad5195ac",
   738 => x"2d720981",
   739 => x"05537280",
   740 => x"2eb53887",
   741 => x"54729c2a",
   742 => x"73842b54",
   743 => x"5271802e",
   744 => x"83388155",
   745 => x"89722587",
   746 => x"38b71252",
   747 => x"97b204b0",
   748 => x"12527480",
   749 => x"2e863871",
   750 => x"5195ac2d",
   751 => x"ff145473",
   752 => x"8025d238",
   753 => x"97cc04b0",
   754 => x"5195ac2d",
   755 => x"800bb3e0",
   756 => x"0c029405",
   757 => x"0d0402c0",
   758 => x"050d0280",
   759 => x"c4055780",
   760 => x"70787084",
   761 => x"055a0872",
   762 => x"415f5d58",
   763 => x"7c708405",
   764 => x"5e085a80",
   765 => x"5b79982a",
   766 => x"7a882b5b",
   767 => x"56758638",
   768 => x"775f99ce",
   769 => x"047d802e",
   770 => x"81a23880",
   771 => x"5e7580e4",
   772 => x"2e8a3875",
   773 => x"80f82e09",
   774 => x"81068938",
   775 => x"76841871",
   776 => x"085e5854",
   777 => x"7580e42e",
   778 => x"9f387580",
   779 => x"e4268a38",
   780 => x"7580e32e",
   781 => x"be3898fe",
   782 => x"047580f3",
   783 => x"2ea33875",
   784 => x"80f82e89",
   785 => x"3898fe04",
   786 => x"8a5398cf",
   787 => x"049053b4",
   788 => x"c0527b51",
   789 => x"96f72db3",
   790 => x"e008b4c0",
   791 => x"5a55998e",
   792 => x"04768418",
   793 => x"71087054",
   794 => x"5b585495",
   795 => x"ce2d8055",
   796 => x"998e0476",
   797 => x"84187108",
   798 => x"58585499",
   799 => x"b904a551",
   800 => x"95ac2d75",
   801 => x"5195ac2d",
   802 => x"82185899",
   803 => x"c10474ff",
   804 => x"16565480",
   805 => x"7425aa38",
   806 => x"78708105",
   807 => x"5a80f52d",
   808 => x"70525695",
   809 => x"ac2d8118",
   810 => x"58998e04",
   811 => x"75a52e09",
   812 => x"81068638",
   813 => x"815e99c1",
   814 => x"04755195",
   815 => x"ac2d8118",
   816 => x"58811b5b",
   817 => x"837b25fe",
   818 => x"ac3875fe",
   819 => x"9f387eb3",
   820 => x"e00c0280",
   821 => x"c0050d04",
   822 => x"02ec050d",
   823 => x"76557480",
   824 => x"f52d5170",
   825 => x"802e81f2",
   826 => x"38b58408",
   827 => x"70828080",
   828 => x"29a9dc08",
   829 => x"05b58008",
   830 => x"11515252",
   831 => x"718f24de",
   832 => x"38747081",
   833 => x"055680f5",
   834 => x"2d527180",
   835 => x"2e81cb38",
   836 => x"71882e09",
   837 => x"81069c38",
   838 => x"800bb580",
   839 => x"0825b838",
   840 => x"ff1151a0",
   841 => x"7181b72d",
   842 => x"b58008ff",
   843 => x"05b5800c",
   844 => x"9aff0471",
   845 => x"8a2e0981",
   846 => x"069d38b5",
   847 => x"84088105",
   848 => x"b5840c80",
   849 => x"0bb5800c",
   850 => x"b5840882",
   851 => x"808029a9",
   852 => x"dc080551",
   853 => x"9aff0471",
   854 => x"71708105",
   855 => x"5381b72d",
   856 => x"b5800881",
   857 => x"05b5800c",
   858 => x"b58008a0",
   859 => x"2e098106",
   860 => x"8e38800b",
   861 => x"b5800cb5",
   862 => x"84088105",
   863 => x"b5840c8f",
   864 => x"0bb58408",
   865 => x"2580c738",
   866 => x"a9dc0882",
   867 => x"80801171",
   868 => x"53555381",
   869 => x"ff527370",
   870 => x"84055508",
   871 => x"71708405",
   872 => x"530cff12",
   873 => x"52718025",
   874 => x"ed388880",
   875 => x"13518f52",
   876 => x"80717084",
   877 => x"05530cff",
   878 => x"12527180",
   879 => x"25f23880",
   880 => x"0bb5800c",
   881 => x"8f0bb584",
   882 => x"0c9e8080",
   883 => x"13518f0b",
   884 => x"b5840825",
   885 => x"feab3899",
   886 => x"de040294",
   887 => x"050d0402",
   888 => x"f4050d02",
   889 => x"930580f5",
   890 => x"2d028c05",
   891 => x"81b72d80",
   892 => x"02840589",
   893 => x"0581b72d",
   894 => x"028c05fc",
   895 => x"055199d8",
   896 => x"2d810bb3",
   897 => x"e00c028c",
   898 => x"050d0402",
   899 => x"fc050d72",
   900 => x"5199d82d",
   901 => x"800bb3e0",
   902 => x"0c028405",
   903 => x"0d0402f8",
   904 => x"050da9dc",
   905 => x"08528ffc",
   906 => x"51807270",
   907 => x"8405540c",
   908 => x"fc115170",
   909 => x"8025f238",
   910 => x"0288050d",
   911 => x"0402fc05",
   912 => x"0d725180",
   913 => x"710c800b",
   914 => x"84120c80",
   915 => x"0b88120c",
   916 => x"800b8c12",
   917 => x"0c028405",
   918 => x"0d0402f0",
   919 => x"050d7570",
   920 => x"08841208",
   921 => x"535353ff",
   922 => x"5471712e",
   923 => x"9b388413",
   924 => x"08708429",
   925 => x"14931180",
   926 => x"f52d8416",
   927 => x"08811187",
   928 => x"0684180c",
   929 => x"52565151",
   930 => x"73b3e00c",
   931 => x"0290050d",
   932 => x"0402f405",
   933 => x"0d747008",
   934 => x"84120853",
   935 => x"53537072",
   936 => x"248f3872",
   937 => x"08841408",
   938 => x"71713152",
   939 => x"52529dbe",
   940 => x"04720884",
   941 => x"14087171",
   942 => x"31880552",
   943 => x"525271b3",
   944 => x"e00c028c",
   945 => x"050d0402",
   946 => x"f8050da2",
   947 => x"ab2da29e",
   948 => x"2de00870",
   949 => x"8b2a7081",
   950 => x"06515252",
   951 => x"70802e9d",
   952 => x"38b9e808",
   953 => x"708429b9",
   954 => x"f8057381",
   955 => x"ff06710c",
   956 => x"5151b9e8",
   957 => x"08811187",
   958 => x"06b9e80c",
   959 => x"51718a2a",
   960 => x"70810651",
   961 => x"5170802e",
   962 => x"a838b9f0",
   963 => x"08b9f408",
   964 => x"52527171",
   965 => x"2e9b38b9",
   966 => x"f0087084",
   967 => x"29ba9805",
   968 => x"7008e00c",
   969 => x"5151b9f0",
   970 => x"08811187",
   971 => x"06b9f00c",
   972 => x"51a2a52d",
   973 => x"0288050d",
   974 => x"0402f405",
   975 => x"0d74538c",
   976 => x"13088111",
   977 => x"87068815",
   978 => x"08545151",
   979 => x"71712eef",
   980 => x"38a2ab2d",
   981 => x"8c130870",
   982 => x"84291477",
   983 => x"b0120c51",
   984 => x"518c1308",
   985 => x"81118706",
   986 => x"8c150c51",
   987 => x"9dc72da2",
   988 => x"a52d028c",
   989 => x"050d0402",
   990 => x"fc050db9",
   991 => x"e8519cbd",
   992 => x"2d9dc751",
   993 => x"a29a2da1",
   994 => x"d22d0284",
   995 => x"050d0402",
   996 => x"e4050d80",
   997 => x"57a19d04",
   998 => x"b3e00881",
   999 => x"f02e0981",
  1000 => x"06893881",
  1001 => x"0bb5900c",
  1002 => x"a19d04b3",
  1003 => x"e00881e0",
  1004 => x"2e098106",
  1005 => x"8938810b",
  1006 => x"b5940ca1",
  1007 => x"9d04b3e0",
  1008 => x"0854b594",
  1009 => x"08802e88",
  1010 => x"38b3e008",
  1011 => x"81800554",
  1012 => x"b5900881",
  1013 => x"9c38830b",
  1014 => x"a9e01581",
  1015 => x"b72d7480",
  1016 => x"ff24b138",
  1017 => x"b58c0882",
  1018 => x"2a708106",
  1019 => x"b5880870",
  1020 => x"872b8180",
  1021 => x"07781182",
  1022 => x"2b515658",
  1023 => x"5154738b",
  1024 => x"38758180",
  1025 => x"29157082",
  1026 => x"2b5153ab",
  1027 => x"e0130853",
  1028 => x"7281b638",
  1029 => x"800bb594",
  1030 => x"0c7480d9",
  1031 => x"2e80c738",
  1032 => x"7480d924",
  1033 => x"8f387492",
  1034 => x"2ebc3874",
  1035 => x"80d82e93",
  1036 => x"38a19804",
  1037 => x"7480f72e",
  1038 => x"a0387480",
  1039 => x"fe2e8f38",
  1040 => x"a19804b5",
  1041 => x"8c088432",
  1042 => x"b58c0ca0",
  1043 => x"e104b58c",
  1044 => x"088132b5",
  1045 => x"8c0ca0e1",
  1046 => x"04b58c08",
  1047 => x"8232b58c",
  1048 => x"0c8157a1",
  1049 => x"9804b588",
  1050 => x"088107b5",
  1051 => x"880ca198",
  1052 => x"04a9e014",
  1053 => x"80f52d81",
  1054 => x"fe065372",
  1055 => x"a9e01581",
  1056 => x"b72d7492",
  1057 => x"2e8a3874",
  1058 => x"80d92e09",
  1059 => x"81068938",
  1060 => x"b58808fe",
  1061 => x"06b5880c",
  1062 => x"800bb590",
  1063 => x"0cb9e851",
  1064 => x"9cda2db3",
  1065 => x"e00855b3",
  1066 => x"e008ff24",
  1067 => x"fdea3876",
  1068 => x"802e9438",
  1069 => x"81ed52b9",
  1070 => x"e8519eb9",
  1071 => x"2db58c08",
  1072 => x"52b9e851",
  1073 => x"9eb92d80",
  1074 => x"5372b3e0",
  1075 => x"0c029c05",
  1076 => x"0d0402fc",
  1077 => x"050d8051",
  1078 => x"800ba9e0",
  1079 => x"1281b72d",
  1080 => x"81115181",
  1081 => x"ff7125f0",
  1082 => x"38028405",
  1083 => x"0d0402f4",
  1084 => x"050d7451",
  1085 => x"a2ab2da9",
  1086 => x"e01180f5",
  1087 => x"2d7081ff",
  1088 => x"0671fd06",
  1089 => x"52545271",
  1090 => x"a9e01281",
  1091 => x"b72da2a5",
  1092 => x"2d72b3e0",
  1093 => x"0c028c05",
  1094 => x"0d047198",
  1095 => x"0c04ffb0",
  1096 => x"08b3e00c",
  1097 => x"04810bff",
  1098 => x"b00c0480",
  1099 => x"0bffb00c",
  1100 => x"0402e805",
  1101 => x"0d787871",
  1102 => x"54575372",
  1103 => x"80258438",
  1104 => x"83135271",
  1105 => x"822cff05",
  1106 => x"5372ff2e",
  1107 => x"80c03875",
  1108 => x"70840557",
  1109 => x"08548755",
  1110 => x"739c2ab0",
  1111 => x"0552b972",
  1112 => x"27843887",
  1113 => x"12527151",
  1114 => x"95ac2d73",
  1115 => x"842bff16",
  1116 => x"56547480",
  1117 => x"25e238a0",
  1118 => x"5195ac2d",
  1119 => x"72870652",
  1120 => x"7186388a",
  1121 => x"5195ac2d",
  1122 => x"ff1353a2",
  1123 => x"c9048a51",
  1124 => x"95ac2d02",
  1125 => x"98050d04",
  1126 => x"b3ec0802",
  1127 => x"b3ec0cff",
  1128 => x"3d0d800b",
  1129 => x"b3ec08fc",
  1130 => x"050cb3ec",
  1131 => x"08880508",
  1132 => x"8106ff11",
  1133 => x"700970b3",
  1134 => x"ec088c05",
  1135 => x"0806b3ec",
  1136 => x"08fc0508",
  1137 => x"11b3ec08",
  1138 => x"fc050cb3",
  1139 => x"ec088805",
  1140 => x"08812ab3",
  1141 => x"ec088805",
  1142 => x"0cb3ec08",
  1143 => x"8c050810",
  1144 => x"b3ec088c",
  1145 => x"050c5151",
  1146 => x"5151b3ec",
  1147 => x"08880508",
  1148 => x"802e8438",
  1149 => x"ffb439b3",
  1150 => x"ec08fc05",
  1151 => x"0870b3e0",
  1152 => x"0c51833d",
  1153 => x"0db3ec0c",
  1154 => x"04000000",
  1155 => x"00ffffff",
  1156 => x"ff00ffff",
  1157 => x"ffff00ff",
  1158 => x"ffffff00",
  1159 => x"496e6974",
  1160 => x"69616c69",
  1161 => x"73696e67",
  1162 => x"2050532f",
  1163 => x"3220696e",
  1164 => x"74657266",
  1165 => x"6163652e",
  1166 => x"2e2e0a00",
  1167 => x"496e6974",
  1168 => x"69616c69",
  1169 => x"7a696e67",
  1170 => x"20534420",
  1171 => x"63617264",
  1172 => x"0a000000",
  1173 => x"48756e74",
  1174 => x"696e6720",
  1175 => x"666f7220",
  1176 => x"70617274",
  1177 => x"6974696f",
  1178 => x"6e0a0000",
  1179 => x"42494f53",
  1180 => x"5041434b",
  1181 => x"524f4d00",
  1182 => x"4f70656e",
  1183 => x"65642066",
  1184 => x"696c652c",
  1185 => x"206c6f61",
  1186 => x"64696e67",
  1187 => x"2e2e2e0a",
  1188 => x"00000000",
  1189 => x"52656164",
  1190 => x"20626c6f",
  1191 => x"636b2066",
  1192 => x"61696c65",
  1193 => x"640a0000",
  1194 => x"4c6f6164",
  1195 => x"696e6720",
  1196 => x"42494f53",
  1197 => x"20666169",
  1198 => x"6c65640a",
  1199 => x"00000000",
  1200 => x"52656164",
  1201 => x"696e6720",
  1202 => x"4d42520a",
  1203 => x"00000000",
  1204 => x"52656164",
  1205 => x"206f6620",
  1206 => x"4d425220",
  1207 => x"6661696c",
  1208 => x"65640a00",
  1209 => x"4d425220",
  1210 => x"73756363",
  1211 => x"65737366",
  1212 => x"756c6c79",
  1213 => x"20726561",
  1214 => x"640a0000",
  1215 => x"46415431",
  1216 => x"36202020",
  1217 => x"00000000",
  1218 => x"46415433",
  1219 => x"32202020",
  1220 => x"00000000",
  1221 => x"50617274",
  1222 => x"6974696f",
  1223 => x"6e636f75",
  1224 => x"6e742025",
  1225 => x"640a0000",
  1226 => x"4e6f2070",
  1227 => x"61727469",
  1228 => x"74696f6e",
  1229 => x"20736967",
  1230 => x"6e617475",
  1231 => x"72652066",
  1232 => x"6f756e64",
  1233 => x"0a000000",
  1234 => x"52656164",
  1235 => x"696e6720",
  1236 => x"626f6f74",
  1237 => x"20736563",
  1238 => x"746f7220",
  1239 => x"25640a00",
  1240 => x"52656164",
  1241 => x"20626f6f",
  1242 => x"74207365",
  1243 => x"63746f72",
  1244 => x"2066726f",
  1245 => x"6d206669",
  1246 => x"72737420",
  1247 => x"70617274",
  1248 => x"6974696f",
  1249 => x"6e0a0000",
  1250 => x"48756e74",
  1251 => x"696e6720",
  1252 => x"666f7220",
  1253 => x"66696c65",
  1254 => x"73797374",
  1255 => x"656d0a00",
  1256 => x"556e7375",
  1257 => x"70706f72",
  1258 => x"74656420",
  1259 => x"70617274",
  1260 => x"6974696f",
  1261 => x"6e207479",
  1262 => x"7065210d",
  1263 => x"00000000",
  1264 => x"436c7573",
  1265 => x"74657220",
  1266 => x"73697a65",
  1267 => x"3a202564",
  1268 => x"2c20436c",
  1269 => x"75737465",
  1270 => x"72206d61",
  1271 => x"736b2c20",
  1272 => x"25640a00",
  1273 => x"47657443",
  1274 => x"6c757374",
  1275 => x"65722072",
  1276 => x"65616469",
  1277 => x"6e672073",
  1278 => x"6563746f",
  1279 => x"72202564",
  1280 => x"0a000000",
  1281 => x"52656164",
  1282 => x"696e6720",
  1283 => x"64697265",
  1284 => x"63746f72",
  1285 => x"79207365",
  1286 => x"63746f72",
  1287 => x"2025640a",
  1288 => x"00000000",
  1289 => x"47657446",
  1290 => x"41544c69",
  1291 => x"6e6b2072",
  1292 => x"65747572",
  1293 => x"6e656420",
  1294 => x"25640a00",
  1295 => x"436d645f",
  1296 => x"696e6974",
  1297 => x"0a000000",
  1298 => x"636d645f",
  1299 => x"434d4438",
  1300 => x"20726573",
  1301 => x"706f6e73",
  1302 => x"653a2025",
  1303 => x"640a0000",
  1304 => x"434d4438",
  1305 => x"5f342072",
  1306 => x"6573706f",
  1307 => x"6e73653a",
  1308 => x"2025640a",
  1309 => x"00000000",
  1310 => x"53444843",
  1311 => x"20496e69",
  1312 => x"7469616c",
  1313 => x"697a6174",
  1314 => x"696f6e20",
  1315 => x"6572726f",
  1316 => x"72210a00",
  1317 => x"434d4435",
  1318 => x"38202564",
  1319 => x"0a202000",
  1320 => x"434d4435",
  1321 => x"385f3220",
  1322 => x"25640a20",
  1323 => x"20000000",
  1324 => x"53504920",
  1325 => x"496e6974",
  1326 => x"28290a00",
  1327 => x"52656164",
  1328 => x"20636f6d",
  1329 => x"6d616e64",
  1330 => x"20666169",
  1331 => x"6c656420",
  1332 => x"61742025",
  1333 => x"64202825",
  1334 => x"64290a00",
  1335 => x"ffffe000",
  1336 => x"00000000",
  1337 => x"00000000",
  1338 => x"00000000",
  1339 => x"00000000",
  1340 => x"00000000",
  1341 => x"00000000",
  1342 => x"00000000",
  1343 => x"00000000",
  1344 => x"00000000",
  1345 => x"00000000",
  1346 => x"00000000",
  1347 => x"00000000",
  1348 => x"00000000",
  1349 => x"00000000",
  1350 => x"00000000",
  1351 => x"00000000",
  1352 => x"00000000",
  1353 => x"00000000",
  1354 => x"00000000",
  1355 => x"00000000",
  1356 => x"00000000",
  1357 => x"00000000",
  1358 => x"00000000",
  1359 => x"00000000",
  1360 => x"00000000",
  1361 => x"00000000",
  1362 => x"00000000",
  1363 => x"00000000",
  1364 => x"00000000",
  1365 => x"00000000",
  1366 => x"00000000",
  1367 => x"00000000",
  1368 => x"00000000",
  1369 => x"00000000",
  1370 => x"00000000",
  1371 => x"00000000",
  1372 => x"00000000",
  1373 => x"00000000",
  1374 => x"00000000",
  1375 => x"00000000",
  1376 => x"00000000",
  1377 => x"00000000",
  1378 => x"00000000",
  1379 => x"00000000",
  1380 => x"00000000",
  1381 => x"00000000",
  1382 => x"00000000",
  1383 => x"00000000",
  1384 => x"00000000",
  1385 => x"00000000",
  1386 => x"00000000",
  1387 => x"00000000",
  1388 => x"00000000",
  1389 => x"00000000",
  1390 => x"00000000",
  1391 => x"00000000",
  1392 => x"00000000",
  1393 => x"00000000",
  1394 => x"00000000",
  1395 => x"00000000",
  1396 => x"00000000",
  1397 => x"00000000",
  1398 => x"00000000",
  1399 => x"00000000",
  1400 => x"00000000",
  1401 => x"00000000",
  1402 => x"00000000",
  1403 => x"00000000",
  1404 => x"00000000",
  1405 => x"00000000",
  1406 => x"00000000",
  1407 => x"00000000",
  1408 => x"00000000",
  1409 => x"00000000",
  1410 => x"00000000",
  1411 => x"00000000",
  1412 => x"00000000",
  1413 => x"00000009",
  1414 => x"00000000",
  1415 => x"00000000",
  1416 => x"00000000",
  1417 => x"00000000",
  1418 => x"00000000",
  1419 => x"00000000",
  1420 => x"00000000",
  1421 => x"00000071",
  1422 => x"00000031",
  1423 => x"00000000",
  1424 => x"00000000",
  1425 => x"00000000",
  1426 => x"0000007a",
  1427 => x"00000073",
  1428 => x"00000061",
  1429 => x"00000077",
  1430 => x"00000032",
  1431 => x"00000000",
  1432 => x"00000000",
  1433 => x"00000063",
  1434 => x"00000078",
  1435 => x"00000064",
  1436 => x"00000065",
  1437 => x"00000034",
  1438 => x"00000033",
  1439 => x"00000000",
  1440 => x"00000000",
  1441 => x"00000020",
  1442 => x"00000076",
  1443 => x"00000066",
  1444 => x"00000074",
  1445 => x"00000072",
  1446 => x"00000035",
  1447 => x"00000000",
  1448 => x"00000000",
  1449 => x"0000006e",
  1450 => x"00000062",
  1451 => x"00000068",
  1452 => x"00000067",
  1453 => x"00000079",
  1454 => x"00000036",
  1455 => x"00000000",
  1456 => x"00000000",
  1457 => x"00000000",
  1458 => x"0000006d",
  1459 => x"0000006a",
  1460 => x"00000075",
  1461 => x"00000037",
  1462 => x"00000038",
  1463 => x"00000000",
  1464 => x"00000000",
  1465 => x"0000002c",
  1466 => x"0000006b",
  1467 => x"00000069",
  1468 => x"0000006f",
  1469 => x"00000030",
  1470 => x"00000039",
  1471 => x"00000000",
  1472 => x"00000000",
  1473 => x"0000002e",
  1474 => x"0000002f",
  1475 => x"0000006c",
  1476 => x"0000003b",
  1477 => x"00000070",
  1478 => x"0000002d",
  1479 => x"00000000",
  1480 => x"00000000",
  1481 => x"00000000",
  1482 => x"00000027",
  1483 => x"00000000",
  1484 => x"0000005b",
  1485 => x"0000003d",
  1486 => x"00000000",
  1487 => x"00000000",
  1488 => x"00000000",
  1489 => x"00000000",
  1490 => x"0000000a",
  1491 => x"0000005d",
  1492 => x"00000000",
  1493 => x"00000023",
  1494 => x"00000000",
  1495 => x"00000000",
  1496 => x"00000000",
  1497 => x"00000000",
  1498 => x"00000000",
  1499 => x"00000000",
  1500 => x"00000000",
  1501 => x"00000000",
  1502 => x"00000008",
  1503 => x"00000000",
  1504 => x"00000000",
  1505 => x"00000031",
  1506 => x"00000000",
  1507 => x"00000034",
  1508 => x"00000037",
  1509 => x"00000000",
  1510 => x"00000000",
  1511 => x"00000000",
  1512 => x"00000030",
  1513 => x"0000002e",
  1514 => x"00000032",
  1515 => x"00000035",
  1516 => x"00000036",
  1517 => x"00000038",
  1518 => x"0000001b",
  1519 => x"00000000",
  1520 => x"00000000",
  1521 => x"0000002b",
  1522 => x"00000033",
  1523 => x"00000000",
  1524 => x"0000002a",
  1525 => x"00000039",
  1526 => x"00000000",
  1527 => x"00000000",
  1528 => x"00000000",
  1529 => x"00000000",
  1530 => x"00000000",
  1531 => x"00000000",
  1532 => x"00000000",
  1533 => x"00000000",
  1534 => x"00000000",
  1535 => x"00000000",
  1536 => x"00000000",
  1537 => x"00000000",
  1538 => x"00000000",
  1539 => x"00000000",
  1540 => x"00000000",
  1541 => x"00000008",
  1542 => x"00000000",
  1543 => x"00000000",
  1544 => x"00000000",
  1545 => x"00000000",
  1546 => x"00000000",
  1547 => x"00000000",
  1548 => x"00000000",
  1549 => x"00000051",
  1550 => x"00000021",
  1551 => x"00000000",
  1552 => x"00000000",
  1553 => x"00000000",
  1554 => x"0000005a",
  1555 => x"00000053",
  1556 => x"00000041",
  1557 => x"00000057",
  1558 => x"00000022",
  1559 => x"00000000",
  1560 => x"00000000",
  1561 => x"00000043",
  1562 => x"00000058",
  1563 => x"00000044",
  1564 => x"00000045",
  1565 => x"00000024",
  1566 => x"000000a3",
  1567 => x"00000000",
  1568 => x"00000000",
  1569 => x"00000020",
  1570 => x"00000056",
  1571 => x"00000046",
  1572 => x"00000054",
  1573 => x"00000052",
  1574 => x"00000025",
  1575 => x"00000000",
  1576 => x"00000000",
  1577 => x"0000004e",
  1578 => x"00000042",
  1579 => x"00000048",
  1580 => x"00000047",
  1581 => x"00000059",
  1582 => x"0000005e",
  1583 => x"00000000",
  1584 => x"00000000",
  1585 => x"00000000",
  1586 => x"0000004d",
  1587 => x"0000004a",
  1588 => x"00000055",
  1589 => x"00000026",
  1590 => x"0000002a",
  1591 => x"00000000",
  1592 => x"00000000",
  1593 => x"0000003c",
  1594 => x"0000004b",
  1595 => x"00000049",
  1596 => x"0000004f",
  1597 => x"00000029",
  1598 => x"00000028",
  1599 => x"00000000",
  1600 => x"00000000",
  1601 => x"0000003e",
  1602 => x"0000003f",
  1603 => x"0000004c",
  1604 => x"0000003a",
  1605 => x"00000050",
  1606 => x"0000005f",
  1607 => x"00000000",
  1608 => x"00000000",
  1609 => x"00000000",
  1610 => x"0000003f",
  1611 => x"00000000",
  1612 => x"0000007b",
  1613 => x"0000002b",
  1614 => x"00000000",
  1615 => x"00000000",
  1616 => x"00000000",
  1617 => x"00000000",
  1618 => x"0000000a",
  1619 => x"0000007d",
  1620 => x"00000000",
  1621 => x"0000007e",
  1622 => x"00000000",
  1623 => x"00000000",
  1624 => x"00000000",
  1625 => x"00000000",
  1626 => x"00000000",
  1627 => x"00000000",
  1628 => x"00000000",
  1629 => x"00000000",
  1630 => x"00000009",
  1631 => x"00000000",
  1632 => x"00000000",
  1633 => x"00000031",
  1634 => x"00000000",
  1635 => x"00000034",
  1636 => x"00000037",
  1637 => x"00000000",
  1638 => x"00000000",
  1639 => x"00000000",
  1640 => x"00000030",
  1641 => x"0000002e",
  1642 => x"00000032",
  1643 => x"00000035",
  1644 => x"00000036",
  1645 => x"00000038",
  1646 => x"0000001b",
  1647 => x"00000000",
  1648 => x"00000000",
  1649 => x"0000002b",
  1650 => x"00000033",
  1651 => x"00000000",
  1652 => x"0000002a",
  1653 => x"00000039",
  1654 => x"00000000",
  1655 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

