-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b0bb5",
     9 => x"d0080b0b",
    10 => x"0bb5d408",
    11 => x"0b0b0bb5",
    12 => x"d8080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"b5d80c0b",
    16 => x"0b0bb5d4",
    17 => x"0c0b0b0b",
    18 => x"b5d00c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0babf0",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"b5d070bb",
    57 => x"f0278b38",
    58 => x"80717084",
    59 => x"05530c81",
    60 => x"e2048c51",
    61 => x"8af10402",
    62 => x"fc050df8",
    63 => x"80518f0b",
    64 => x"b5e00c9f",
    65 => x"0bb5e40c",
    66 => x"a0717081",
    67 => x"055334b5",
    68 => x"e408ff05",
    69 => x"b5e40cb5",
    70 => x"e4088025",
    71 => x"eb38b5e0",
    72 => x"08ff05b5",
    73 => x"e00cb5e0",
    74 => x"088025d7",
    75 => x"38028405",
    76 => x"0d0402f0",
    77 => x"050df880",
    78 => x"53f8a054",
    79 => x"83bf5273",
    80 => x"70810555",
    81 => x"33517073",
    82 => x"70810555",
    83 => x"34ff1252",
    84 => x"718025eb",
    85 => x"38fbc053",
    86 => x"9f52a073",
    87 => x"70810555",
    88 => x"34ff1252",
    89 => x"718025f2",
    90 => x"38029005",
    91 => x"0d0402f4",
    92 => x"050d7453",
    93 => x"8e0bb5e0",
    94 => x"08258f38",
    95 => x"82b22db5",
    96 => x"e008ff05",
    97 => x"b5e00c82",
    98 => x"f404b5e0",
    99 => x"08b5e408",
   100 => x"5351728a",
   101 => x"2e098106",
   102 => x"b7387151",
   103 => x"719f24a0",
   104 => x"38b5e008",
   105 => x"a02911f8",
   106 => x"80115151",
   107 => x"a07134b5",
   108 => x"e4088105",
   109 => x"b5e40cb5",
   110 => x"e408519f",
   111 => x"7125e238",
   112 => x"800bb5e4",
   113 => x"0cb5e008",
   114 => x"8105b5e0",
   115 => x"0c83e404",
   116 => x"70a02912",
   117 => x"f8801151",
   118 => x"51727134",
   119 => x"b5e40881",
   120 => x"05b5e40c",
   121 => x"b5e408a0",
   122 => x"2e098106",
   123 => x"8e38800b",
   124 => x"b5e40cb5",
   125 => x"e0088105",
   126 => x"b5e00c02",
   127 => x"8c050d04",
   128 => x"02e8050d",
   129 => x"77795656",
   130 => x"880bfc16",
   131 => x"77712c8f",
   132 => x"06545254",
   133 => x"80537272",
   134 => x"25953871",
   135 => x"53fbe014",
   136 => x"51877134",
   137 => x"8114ff14",
   138 => x"545472f1",
   139 => x"387153f9",
   140 => x"1576712c",
   141 => x"87065351",
   142 => x"71802e8b",
   143 => x"38fbe014",
   144 => x"51717134",
   145 => x"81145472",
   146 => x"8e249538",
   147 => x"8f733153",
   148 => x"fbe01451",
   149 => x"a0713481",
   150 => x"14ff1454",
   151 => x"5472f138",
   152 => x"0298050d",
   153 => x"0402ec05",
   154 => x"0d800bb5",
   155 => x"e80cf68c",
   156 => x"08f69008",
   157 => x"71882c56",
   158 => x"5481ff06",
   159 => x"52737225",
   160 => x"88387154",
   161 => x"820bb5e8",
   162 => x"0c72882c",
   163 => x"7381ff06",
   164 => x"54557473",
   165 => x"258b3872",
   166 => x"b5e80884",
   167 => x"07b5e80c",
   168 => x"5573842b",
   169 => x"86a07125",
   170 => x"83713170",
   171 => x"0b0b0bb3",
   172 => x"900c8171",
   173 => x"2bff05f6",
   174 => x"880cfecc",
   175 => x"13ff122c",
   176 => x"788829ff",
   177 => x"94057081",
   178 => x"2cb5e808",
   179 => x"52585255",
   180 => x"51525476",
   181 => x"802e8538",
   182 => x"70810751",
   183 => x"70f6940c",
   184 => x"71098105",
   185 => x"f6800c72",
   186 => x"098105f6",
   187 => x"840c0294",
   188 => x"050d0402",
   189 => x"f4050d74",
   190 => x"53727081",
   191 => x"055480f5",
   192 => x"2d527180",
   193 => x"2e893871",
   194 => x"5182ee2d",
   195 => x"85f90402",
   196 => x"8c050d04",
   197 => x"02f8050d",
   198 => x"a5c92d80",
   199 => x"da51a780",
   200 => x"2db5d008",
   201 => x"812a7081",
   202 => x"06515271",
   203 => x"802ee938",
   204 => x"0288050d",
   205 => x"0402f405",
   206 => x"0dbbe008",
   207 => x"99c406b4",
   208 => x"ac0b80f5",
   209 => x"2d525270",
   210 => x"802e8638",
   211 => x"71848007",
   212 => x"52b3e40b",
   213 => x"80f52d72",
   214 => x"07b3fc0b",
   215 => x"80f52d70",
   216 => x"812a7081",
   217 => x"06515354",
   218 => x"5270802e",
   219 => x"86387182",
   220 => x"80075272",
   221 => x"81065170",
   222 => x"802e8538",
   223 => x"71880752",
   224 => x"b4880b80",
   225 => x"f52d7084",
   226 => x"2b730781",
   227 => x"8432b5d0",
   228 => x"0c51028c",
   229 => x"050d0402",
   230 => x"f4050d74",
   231 => x"70818432",
   232 => x"bbe00c70",
   233 => x"83065253",
   234 => x"70b3dc0b",
   235 => x"880581b7",
   236 => x"2d72892a",
   237 => x"70810651",
   238 => x"5170b4ac",
   239 => x"0b81b72d",
   240 => x"72832a81",
   241 => x"0673882a",
   242 => x"70810651",
   243 => x"52527080",
   244 => x"2e853871",
   245 => x"82075271",
   246 => x"b3fc0b81",
   247 => x"b72d7284",
   248 => x"2c708306",
   249 => x"515170b4",
   250 => x"880b81b7",
   251 => x"2d70b5d0",
   252 => x"0c028c05",
   253 => x"0d0402d4",
   254 => x"050daed4",
   255 => x"5185f32d",
   256 => x"9b852db5",
   257 => x"d008802e",
   258 => x"82ab3886",
   259 => x"b52db5d0",
   260 => x"08538de0",
   261 => x"2db5d008",
   262 => x"54b5d008",
   263 => x"802e8297",
   264 => x"389dc82d",
   265 => x"b5d00880",
   266 => x"2e8738ae",
   267 => x"ec5188be",
   268 => x"0496e72d",
   269 => x"b5d00880",
   270 => x"2e9c38af",
   271 => x"ac5185f3",
   272 => x"2d86942d",
   273 => x"72840753",
   274 => x"810bfec4",
   275 => x"0c72fec0",
   276 => x"0c725187",
   277 => x"972d840b",
   278 => x"fec40caf",
   279 => x"f45185f3",
   280 => x"2db08c52",
   281 => x"b5f05193",
   282 => x"fc2db5d0",
   283 => x"089838b0",
   284 => x"985185f3",
   285 => x"2db0b052",
   286 => x"b5f05193",
   287 => x"fc2db5d0",
   288 => x"08802e81",
   289 => x"b038b0bc",
   290 => x"5185f32d",
   291 => x"b5f40857",
   292 => x"8077595a",
   293 => x"767a2e8b",
   294 => x"38811a78",
   295 => x"812a595a",
   296 => x"77f738f7",
   297 => x"1a5a8077",
   298 => x"25818038",
   299 => x"79527751",
   300 => x"84802db5",
   301 => x"fc52b5f0",
   302 => x"5196c12d",
   303 => x"b5d00853",
   304 => x"b5d00880",
   305 => x"2e80c938",
   306 => x"b5fc5b80",
   307 => x"5989fd04",
   308 => x"7a708405",
   309 => x"5c087081",
   310 => x"ff067188",
   311 => x"2c7081ff",
   312 => x"0673902c",
   313 => x"7081ff06",
   314 => x"75982afe",
   315 => x"c80cfec8",
   316 => x"0c58fec8",
   317 => x"0c57fec8",
   318 => x"0c841a5a",
   319 => x"53765384",
   320 => x"80772584",
   321 => x"38848053",
   322 => x"727924c4",
   323 => x"388a9b04",
   324 => x"b0d85185",
   325 => x"f32d7254",
   326 => x"8ab704b5",
   327 => x"f0519694",
   328 => x"2dfc8017",
   329 => x"81195957",
   330 => x"89a60482",
   331 => x"0bfec40c",
   332 => x"81548ab7",
   333 => x"04805473",
   334 => x"b5d00c02",
   335 => x"ac050d04",
   336 => x"02f8050d",
   337 => x"a7d02d81",
   338 => x"f72d8151",
   339 => x"84e52dfe",
   340 => x"c4528172",
   341 => x"0ca58d2d",
   342 => x"a58d2d84",
   343 => x"720c87f6",
   344 => x"2db39451",
   345 => x"a8e92d80",
   346 => x"5184e52d",
   347 => x"0288050d",
   348 => x"0402ec05",
   349 => x"0d8cb851",
   350 => x"87972d81",
   351 => x"0bfec40c",
   352 => x"8cb80bfe",
   353 => x"c00c840b",
   354 => x"fec40c83",
   355 => x"0bfecc0c",
   356 => x"a5a82da7",
   357 => x"c42da58d",
   358 => x"2da58d2d",
   359 => x"81f72d81",
   360 => x"5184e52d",
   361 => x"a58d2da5",
   362 => x"8d2d8151",
   363 => x"84e52d87",
   364 => x"f62db5d0",
   365 => x"08802e81",
   366 => x"d4388051",
   367 => x"84e52db3",
   368 => x"9451a8e9",
   369 => x"2dbbc808",
   370 => x"09708306",
   371 => x"fecc0c52",
   372 => x"bbc00889",
   373 => x"38bbc408",
   374 => x"802e80e2",
   375 => x"38fed008",
   376 => x"70810651",
   377 => x"5271802e",
   378 => x"80d438a7",
   379 => x"ca2dbbc0",
   380 => x"0870bbc4",
   381 => x"08705755",
   382 => x"565280ff",
   383 => x"72258438",
   384 => x"80ff5280",
   385 => x"ff732584",
   386 => x"3880ff53",
   387 => x"71ff8025",
   388 => x"8438ff80",
   389 => x"5272ff80",
   390 => x"258438ff",
   391 => x"80537472",
   392 => x"31bbc00c",
   393 => x"737331bb",
   394 => x"c40ca7c4",
   395 => x"2d71882b",
   396 => x"83fe8006",
   397 => x"7381ff06",
   398 => x"7107fed0",
   399 => x"0c52a5c9",
   400 => x"2da8f92d",
   401 => x"b5d00853",
   402 => x"86b52db5",
   403 => x"d008fec0",
   404 => x"0c86b52d",
   405 => x"b5d008b5",
   406 => x"ec082e9c",
   407 => x"38b5d008",
   408 => x"b5ec0c84",
   409 => x"52725184",
   410 => x"e52da58d",
   411 => x"2da58d2d",
   412 => x"ff125271",
   413 => x"8025ee38",
   414 => x"72802e89",
   415 => x"388a0bfe",
   416 => x"c40c8bc5",
   417 => x"04820bfe",
   418 => x"c40c8bc5",
   419 => x"04b0ec51",
   420 => x"85f32d82",
   421 => x"0bfec40c",
   422 => x"800bb5d0",
   423 => x"0c029405",
   424 => x"0d0402e8",
   425 => x"050d7779",
   426 => x"7b585555",
   427 => x"80537276",
   428 => x"25a33874",
   429 => x"70810556",
   430 => x"80f52d74",
   431 => x"70810556",
   432 => x"80f52d52",
   433 => x"5271712e",
   434 => x"86388151",
   435 => x"8dd70481",
   436 => x"13538dae",
   437 => x"04805170",
   438 => x"b5d00c02",
   439 => x"98050d04",
   440 => x"02d8050d",
   441 => x"800bba84",
   442 => x"0cb5fc52",
   443 => x"80519ca5",
   444 => x"2db5d008",
   445 => x"54b5d008",
   446 => x"8c38b184",
   447 => x"5185f32d",
   448 => x"73559385",
   449 => x"04805681",
   450 => x"0bbaa80c",
   451 => x"8853b198",
   452 => x"52b6b251",
   453 => x"8da22db5",
   454 => x"d008762e",
   455 => x"09810687",
   456 => x"38b5d008",
   457 => x"baa80c88",
   458 => x"53b1a452",
   459 => x"b6ce518d",
   460 => x"a22db5d0",
   461 => x"088738b5",
   462 => x"d008baa8",
   463 => x"0cbaa808",
   464 => x"52b1b051",
   465 => x"9fc22dba",
   466 => x"a808802e",
   467 => x"80f638b9",
   468 => x"c20b80f5",
   469 => x"2db9c30b",
   470 => x"80f52d71",
   471 => x"982b7190",
   472 => x"2b07b9c4",
   473 => x"0b80f52d",
   474 => x"70882b72",
   475 => x"07b9c50b",
   476 => x"80f52d71",
   477 => x"07b9fa0b",
   478 => x"80f52db9",
   479 => x"fb0b80f5",
   480 => x"2d71882b",
   481 => x"07535f54",
   482 => x"525a5657",
   483 => x"557381ab",
   484 => x"aa2e0981",
   485 => x"068d3875",
   486 => x"519e972d",
   487 => x"b5d00856",
   488 => x"8fb00473",
   489 => x"82d4d52e",
   490 => x"8738b1c8",
   491 => x"518ff104",
   492 => x"b5fc5275",
   493 => x"519ca52d",
   494 => x"b5d00855",
   495 => x"b5d00880",
   496 => x"2e83c238",
   497 => x"8853b1a4",
   498 => x"52b6ce51",
   499 => x"8da22db5",
   500 => x"d0088938",
   501 => x"810bba84",
   502 => x"0c8ff704",
   503 => x"8853b198",
   504 => x"52b6b251",
   505 => x"8da22db5",
   506 => x"d008802e",
   507 => x"8a38b1e8",
   508 => x"5185f32d",
   509 => x"90d104b9",
   510 => x"fa0b80f5",
   511 => x"2d547380",
   512 => x"d52e0981",
   513 => x"0680ca38",
   514 => x"b9fb0b80",
   515 => x"f52d5473",
   516 => x"81aa2e09",
   517 => x"8106ba38",
   518 => x"800bb5fc",
   519 => x"0b80f52d",
   520 => x"56547481",
   521 => x"e92e8338",
   522 => x"81547481",
   523 => x"eb2e8c38",
   524 => x"80557375",
   525 => x"2e098106",
   526 => x"82cb38b6",
   527 => x"870b80f5",
   528 => x"2d55748d",
   529 => x"38b6880b",
   530 => x"80f52d54",
   531 => x"73822e86",
   532 => x"38805593",
   533 => x"8504b689",
   534 => x"0b80f52d",
   535 => x"70b9fc0c",
   536 => x"ff05ba80",
   537 => x"0cb68a0b",
   538 => x"80f52db6",
   539 => x"8b0b80f5",
   540 => x"2d587605",
   541 => x"77828029",
   542 => x"0570ba88",
   543 => x"0cb68c0b",
   544 => x"80f52d70",
   545 => x"ba9c0cba",
   546 => x"84085957",
   547 => x"5876802e",
   548 => x"81a33888",
   549 => x"53b1a452",
   550 => x"b6ce518d",
   551 => x"a22db5d0",
   552 => x"0881e238",
   553 => x"b9fc0870",
   554 => x"842bbaa0",
   555 => x"0c70ba98",
   556 => x"0cb6a10b",
   557 => x"80f52db6",
   558 => x"a00b80f5",
   559 => x"2d718280",
   560 => x"2905b6a2",
   561 => x"0b80f52d",
   562 => x"70848080",
   563 => x"2912b6a3",
   564 => x"0b80f52d",
   565 => x"7081800a",
   566 => x"291270ba",
   567 => x"a40cba9c",
   568 => x"087129ba",
   569 => x"88080570",
   570 => x"ba8c0cb6",
   571 => x"a90b80f5",
   572 => x"2db6a80b",
   573 => x"80f52d71",
   574 => x"82802905",
   575 => x"b6aa0b80",
   576 => x"f52d7084",
   577 => x"80802912",
   578 => x"b6ab0b80",
   579 => x"f52d7098",
   580 => x"2b81f00a",
   581 => x"06720570",
   582 => x"ba900cfe",
   583 => x"117e2977",
   584 => x"05ba940c",
   585 => x"52595243",
   586 => x"545e5152",
   587 => x"59525d57",
   588 => x"59579383",
   589 => x"04b68e0b",
   590 => x"80f52db6",
   591 => x"8d0b80f5",
   592 => x"2d718280",
   593 => x"290570ba",
   594 => x"a00c70a0",
   595 => x"2983ff05",
   596 => x"70892a70",
   597 => x"ba980cb6",
   598 => x"930b80f5",
   599 => x"2db6920b",
   600 => x"80f52d71",
   601 => x"82802905",
   602 => x"70baa40c",
   603 => x"7b71291e",
   604 => x"70ba940c",
   605 => x"7dba900c",
   606 => x"7305ba8c",
   607 => x"0c555e51",
   608 => x"51555581",
   609 => x"5574b5d0",
   610 => x"0c02a805",
   611 => x"0d0402ec",
   612 => x"050d7670",
   613 => x"872c7180",
   614 => x"ff065556",
   615 => x"54ba8408",
   616 => x"8a387388",
   617 => x"2c7481ff",
   618 => x"065455b5",
   619 => x"fc52ba88",
   620 => x"0815519c",
   621 => x"a52db5d0",
   622 => x"0854b5d0",
   623 => x"08802eb3",
   624 => x"38ba8408",
   625 => x"802e9838",
   626 => x"728429b5",
   627 => x"fc057008",
   628 => x"52539e97",
   629 => x"2db5d008",
   630 => x"f00a0653",
   631 => x"93f10472",
   632 => x"10b5fc05",
   633 => x"7080e02d",
   634 => x"52539ec7",
   635 => x"2db5d008",
   636 => x"53725473",
   637 => x"b5d00c02",
   638 => x"94050d04",
   639 => x"02c8050d",
   640 => x"7f615f5b",
   641 => x"800bba90",
   642 => x"08ba9408",
   643 => x"595d56ba",
   644 => x"8408762e",
   645 => x"8a38b9fc",
   646 => x"08842b58",
   647 => x"94a504ba",
   648 => x"9808842b",
   649 => x"58805978",
   650 => x"782781a9",
   651 => x"38788f06",
   652 => x"a0175754",
   653 => x"738f38b5",
   654 => x"fc527651",
   655 => x"8117579c",
   656 => x"a52db5fc",
   657 => x"56807680",
   658 => x"f52d5654",
   659 => x"74742e83",
   660 => x"38815474",
   661 => x"81e52e80",
   662 => x"f6388170",
   663 => x"7506555d",
   664 => x"73802e80",
   665 => x"ea388b16",
   666 => x"80f52d98",
   667 => x"065a7980",
   668 => x"de388b53",
   669 => x"7d527551",
   670 => x"8da22db5",
   671 => x"d00880cf",
   672 => x"389c1608",
   673 => x"519e972d",
   674 => x"b5d00884",
   675 => x"1c0c9a16",
   676 => x"80e02d51",
   677 => x"9ec72db5",
   678 => x"d008b5d0",
   679 => x"08881d0c",
   680 => x"b5d00855",
   681 => x"55ba8408",
   682 => x"802e9838",
   683 => x"941680e0",
   684 => x"2d519ec7",
   685 => x"2db5d008",
   686 => x"902b83ff",
   687 => x"f00a0670",
   688 => x"16515473",
   689 => x"881c0c79",
   690 => x"7b0c7c54",
   691 => x"968b0481",
   692 => x"195994a7",
   693 => x"04ba8408",
   694 => x"802eae38",
   695 => x"7b51938e",
   696 => x"2db5d008",
   697 => x"b5d00880",
   698 => x"fffffff8",
   699 => x"06555c73",
   700 => x"80ffffff",
   701 => x"f82e9238",
   702 => x"b5d008fe",
   703 => x"05b9fc08",
   704 => x"29ba8c08",
   705 => x"055794a5",
   706 => x"04805473",
   707 => x"b5d00c02",
   708 => x"b8050d04",
   709 => x"02f4050d",
   710 => x"74700881",
   711 => x"05710c70",
   712 => x"08ba8008",
   713 => x"06535371",
   714 => x"8e388813",
   715 => x"0851938e",
   716 => x"2db5d008",
   717 => x"88140c81",
   718 => x"0bb5d00c",
   719 => x"028c050d",
   720 => x"0402f005",
   721 => x"0d758811",
   722 => x"08fe05b9",
   723 => x"fc0829ba",
   724 => x"8c081172",
   725 => x"08ba8008",
   726 => x"06057955",
   727 => x"5354549c",
   728 => x"a52d0290",
   729 => x"050d04ba",
   730 => x"8408b5d0",
   731 => x"0c0402f4",
   732 => x"050dd452",
   733 => x"81ff720c",
   734 => x"71085381",
   735 => x"ff720c72",
   736 => x"882b83fe",
   737 => x"80067208",
   738 => x"7081ff06",
   739 => x"51525381",
   740 => x"ff720c72",
   741 => x"7107882b",
   742 => x"72087081",
   743 => x"ff065152",
   744 => x"5381ff72",
   745 => x"0c727107",
   746 => x"882b7208",
   747 => x"7081ff06",
   748 => x"7207b5d0",
   749 => x"0c525302",
   750 => x"8c050d04",
   751 => x"02f4050d",
   752 => x"74767181",
   753 => x"ff06d40c",
   754 => x"5353baac",
   755 => x"08853871",
   756 => x"892b5271",
   757 => x"982ad40c",
   758 => x"71902a70",
   759 => x"81ff06d4",
   760 => x"0c517188",
   761 => x"2a7081ff",
   762 => x"06d40c51",
   763 => x"7181ff06",
   764 => x"d40c7290",
   765 => x"2a7081ff",
   766 => x"06d40c51",
   767 => x"d4087081",
   768 => x"ff065151",
   769 => x"82b8bf52",
   770 => x"7081ff2e",
   771 => x"09810694",
   772 => x"3881ff0b",
   773 => x"d40cd408",
   774 => x"7081ff06",
   775 => x"ff145451",
   776 => x"5171e538",
   777 => x"70b5d00c",
   778 => x"028c050d",
   779 => x"0402fc05",
   780 => x"0d81c751",
   781 => x"81ff0bd4",
   782 => x"0cff1151",
   783 => x"708025f4",
   784 => x"38028405",
   785 => x"0d0402f0",
   786 => x"050d98ad",
   787 => x"2d8fcf53",
   788 => x"805287fc",
   789 => x"80f75197",
   790 => x"bc2db5d0",
   791 => x"0854b5d0",
   792 => x"08812e09",
   793 => x"8106a338",
   794 => x"81ff0bd4",
   795 => x"0c820a52",
   796 => x"849c80e9",
   797 => x"5197bc2d",
   798 => x"b5d0088b",
   799 => x"3881ff0b",
   800 => x"d40c7353",
   801 => x"99900498",
   802 => x"ad2dff13",
   803 => x"5372c138",
   804 => x"72b5d00c",
   805 => x"0290050d",
   806 => x"0402f405",
   807 => x"0d81ff0b",
   808 => x"d40c9353",
   809 => x"805287fc",
   810 => x"80c15197",
   811 => x"bc2db5d0",
   812 => x"088b3881",
   813 => x"ff0bd40c",
   814 => x"815399c6",
   815 => x"0498ad2d",
   816 => x"ff135372",
   817 => x"df3872b5",
   818 => x"d00c028c",
   819 => x"050d0402",
   820 => x"f0050d98",
   821 => x"ad2d83aa",
   822 => x"52849c80",
   823 => x"c85197bc",
   824 => x"2db5d008",
   825 => x"812e0981",
   826 => x"06923896",
   827 => x"ee2db5d0",
   828 => x"0883ffff",
   829 => x"06537283",
   830 => x"aa2e9738",
   831 => x"99992d9a",
   832 => x"8d048154",
   833 => x"9afc04b2",
   834 => x"885185f3",
   835 => x"2d80549a",
   836 => x"fc0481ff",
   837 => x"0bd40cb1",
   838 => x"5398c62d",
   839 => x"b5d00880",
   840 => x"2e80ca38",
   841 => x"805287fc",
   842 => x"80fa5197",
   843 => x"bc2db5d0",
   844 => x"08b13881",
   845 => x"ff0bd40c",
   846 => x"d4085381",
   847 => x"ff0bd40c",
   848 => x"81ff0bd4",
   849 => x"0c81ff0b",
   850 => x"d40c81ff",
   851 => x"0bd40c72",
   852 => x"862a7081",
   853 => x"06b5d008",
   854 => x"56515372",
   855 => x"802e9d38",
   856 => x"9a8204b5",
   857 => x"d00852b2",
   858 => x"a4519fc2",
   859 => x"2d72822e",
   860 => x"ff9538ff",
   861 => x"135372ff",
   862 => x"a0387254",
   863 => x"73b5d00c",
   864 => x"0290050d",
   865 => x"0402f405",
   866 => x"0d810bba",
   867 => x"ac0cd008",
   868 => x"708f2a70",
   869 => x"81065151",
   870 => x"5372f338",
   871 => x"72d00c98",
   872 => x"ad2db2b0",
   873 => x"5185f32d",
   874 => x"d008708f",
   875 => x"2a708106",
   876 => x"51515372",
   877 => x"f338810b",
   878 => x"d00c80e3",
   879 => x"53805284",
   880 => x"d480c051",
   881 => x"97bc2db5",
   882 => x"d008812e",
   883 => x"9a387282",
   884 => x"2e098106",
   885 => x"8c38b2cc",
   886 => x"5185f32d",
   887 => x"80539c9c",
   888 => x"04ff1353",
   889 => x"72d73899",
   890 => x"cf2db5d0",
   891 => x"08baac0c",
   892 => x"b5d0088b",
   893 => x"38815287",
   894 => x"fc80d051",
   895 => x"97bc2d81",
   896 => x"ff0bd40c",
   897 => x"d008708f",
   898 => x"2a708106",
   899 => x"51515372",
   900 => x"f33872d0",
   901 => x"0c81ff0b",
   902 => x"d40c8153",
   903 => x"72b5d00c",
   904 => x"028c050d",
   905 => x"0402e005",
   906 => x"0d797b57",
   907 => x"57805881",
   908 => x"ff0bd40c",
   909 => x"d008708f",
   910 => x"2a708106",
   911 => x"51515473",
   912 => x"f3388281",
   913 => x"0bd00c81",
   914 => x"ff0bd40c",
   915 => x"765287fc",
   916 => x"80d15197",
   917 => x"bc2d80db",
   918 => x"c6df55b5",
   919 => x"d008802e",
   920 => x"9038b5d0",
   921 => x"08537652",
   922 => x"b2e4519f",
   923 => x"c22d9dbf",
   924 => x"0481ff0b",
   925 => x"d40cd408",
   926 => x"7081ff06",
   927 => x"51547381",
   928 => x"fe2e0981",
   929 => x"069d3880",
   930 => x"ff5496ee",
   931 => x"2db5d008",
   932 => x"76708405",
   933 => x"580cff14",
   934 => x"54738025",
   935 => x"ed388158",
   936 => x"9da904ff",
   937 => x"155574c9",
   938 => x"3881ff0b",
   939 => x"d40cd008",
   940 => x"708f2a70",
   941 => x"81065151",
   942 => x"5473f338",
   943 => x"73d00c77",
   944 => x"b5d00c02",
   945 => x"a0050d04",
   946 => x"baac08b5",
   947 => x"d00c0402",
   948 => x"e8050d80",
   949 => x"78575575",
   950 => x"70840557",
   951 => x"08538054",
   952 => x"72982a73",
   953 => x"882b5452",
   954 => x"71802ea2",
   955 => x"38c00870",
   956 => x"882a7081",
   957 => x"06515151",
   958 => x"70802ef1",
   959 => x"3871c00c",
   960 => x"81158115",
   961 => x"55558374",
   962 => x"25d63871",
   963 => x"ca3874b5",
   964 => x"d00c0298",
   965 => x"050d0402",
   966 => x"f4050d74",
   967 => x"70882a83",
   968 => x"fe800670",
   969 => x"72982a07",
   970 => x"72882b87",
   971 => x"fc808006",
   972 => x"73982b81",
   973 => x"f00a0671",
   974 => x"730707b5",
   975 => x"d00c5651",
   976 => x"5351028c",
   977 => x"050d0402",
   978 => x"f8050d02",
   979 => x"8e0580f5",
   980 => x"2d74882b",
   981 => x"077083ff",
   982 => x"ff06b5d0",
   983 => x"0c510288",
   984 => x"050d0402",
   985 => x"ec050d76",
   986 => x"53805572",
   987 => x"75258b38",
   988 => x"ad5182ee",
   989 => x"2d720981",
   990 => x"05537280",
   991 => x"2eb53887",
   992 => x"54729c2a",
   993 => x"73842b54",
   994 => x"5271802e",
   995 => x"83388155",
   996 => x"89722587",
   997 => x"38b71252",
   998 => x"9f9e04b0",
   999 => x"12527480",
  1000 => x"2e863871",
  1001 => x"5182ee2d",
  1002 => x"ff145473",
  1003 => x"8025d238",
  1004 => x"9fb804b0",
  1005 => x"5182ee2d",
  1006 => x"800bb5d0",
  1007 => x"0c029405",
  1008 => x"0d0402c0",
  1009 => x"050d0280",
  1010 => x"c4055780",
  1011 => x"70787084",
  1012 => x"055a0872",
  1013 => x"415f5d58",
  1014 => x"7c708405",
  1015 => x"5e085a80",
  1016 => x"5b79982a",
  1017 => x"7a882b5b",
  1018 => x"56758638",
  1019 => x"775fa1ba",
  1020 => x"047d802e",
  1021 => x"81a23880",
  1022 => x"5e7580e4",
  1023 => x"2e8a3875",
  1024 => x"80f82e09",
  1025 => x"81068938",
  1026 => x"76841871",
  1027 => x"085e5854",
  1028 => x"7580e42e",
  1029 => x"9f387580",
  1030 => x"e4268a38",
  1031 => x"7580e32e",
  1032 => x"be38a0ea",
  1033 => x"047580f3",
  1034 => x"2ea33875",
  1035 => x"80f82e89",
  1036 => x"38a0ea04",
  1037 => x"8a53a0bb",
  1038 => x"049053ba",
  1039 => x"b0527b51",
  1040 => x"9ee32db5",
  1041 => x"d008bab0",
  1042 => x"5a55a0fa",
  1043 => x"04768418",
  1044 => x"71087054",
  1045 => x"5b58549d",
  1046 => x"cf2d8055",
  1047 => x"a0fa0476",
  1048 => x"84187108",
  1049 => x"585854a1",
  1050 => x"a504a551",
  1051 => x"82ee2d75",
  1052 => x"5182ee2d",
  1053 => x"821858a1",
  1054 => x"ad0474ff",
  1055 => x"16565480",
  1056 => x"7425aa38",
  1057 => x"78708105",
  1058 => x"5a80f52d",
  1059 => x"70525682",
  1060 => x"ee2d8118",
  1061 => x"58a0fa04",
  1062 => x"75a52e09",
  1063 => x"81068638",
  1064 => x"815ea1ad",
  1065 => x"04755182",
  1066 => x"ee2d8118",
  1067 => x"58811b5b",
  1068 => x"837b25fe",
  1069 => x"ac3875fe",
  1070 => x"9f387eb5",
  1071 => x"d00c0280",
  1072 => x"c0050d04",
  1073 => x"02fc050d",
  1074 => x"72518071",
  1075 => x"0c800b84",
  1076 => x"120c0284",
  1077 => x"050d0402",
  1078 => x"f0050d75",
  1079 => x"70088412",
  1080 => x"08535353",
  1081 => x"ff547171",
  1082 => x"2ea838a7",
  1083 => x"ca2d8413",
  1084 => x"08708429",
  1085 => x"14881170",
  1086 => x"087081ff",
  1087 => x"06841808",
  1088 => x"81118706",
  1089 => x"841a0c53",
  1090 => x"51555151",
  1091 => x"51a7c42d",
  1092 => x"715473b5",
  1093 => x"d00c0290",
  1094 => x"050d0402",
  1095 => x"f4050d74",
  1096 => x"53841308",
  1097 => x"81118706",
  1098 => x"74085451",
  1099 => x"5171712e",
  1100 => x"f038a7ca",
  1101 => x"2d841308",
  1102 => x"70842914",
  1103 => x"88117871",
  1104 => x"0c515151",
  1105 => x"84130881",
  1106 => x"11870684",
  1107 => x"150c51a7",
  1108 => x"c42d028c",
  1109 => x"050d0402",
  1110 => x"f0050da7",
  1111 => x"ca2de008",
  1112 => x"e408718b",
  1113 => x"2a708106",
  1114 => x"51535552",
  1115 => x"70802e9d",
  1116 => x"38baf008",
  1117 => x"708429ba",
  1118 => x"f8057381",
  1119 => x"ff06710c",
  1120 => x"5151baf0",
  1121 => x"08811187",
  1122 => x"06baf00c",
  1123 => x"51738b2a",
  1124 => x"70810651",
  1125 => x"5170802e",
  1126 => x"818938b5",
  1127 => x"80088429",
  1128 => x"bbd00574",
  1129 => x"81ff0671",
  1130 => x"0c51b580",
  1131 => x"088105b5",
  1132 => x"800c850b",
  1133 => x"b4fc0cb5",
  1134 => x"8008b4f8",
  1135 => x"082e0981",
  1136 => x"06818638",
  1137 => x"800bb580",
  1138 => x"0cbbd008",
  1139 => x"708306bb",
  1140 => x"c80c7085",
  1141 => x"2a708106",
  1142 => x"bbc40856",
  1143 => x"51525270",
  1144 => x"802e8e38",
  1145 => x"bbd808fe",
  1146 => x"803213bb",
  1147 => x"c40ca3f8",
  1148 => x"04bbd808",
  1149 => x"13bbc40c",
  1150 => x"71842a70",
  1151 => x"8106bbc0",
  1152 => x"08545151",
  1153 => x"70802e90",
  1154 => x"38bbd408",
  1155 => x"81ff3212",
  1156 => x"8105bbc0",
  1157 => x"0ca4c904",
  1158 => x"71bbd408",
  1159 => x"31bbc00c",
  1160 => x"a4c904b4",
  1161 => x"fc08ff05",
  1162 => x"b4fc0cb4",
  1163 => x"fc08ff2e",
  1164 => x"09810695",
  1165 => x"38b58008",
  1166 => x"802e8a38",
  1167 => x"870bb4f8",
  1168 => x"0831b4f8",
  1169 => x"0c70b580",
  1170 => x"0c738a2a",
  1171 => x"70810651",
  1172 => x"5170802e",
  1173 => x"a838bb98",
  1174 => x"08bb9c08",
  1175 => x"52527171",
  1176 => x"2e9b38bb",
  1177 => x"98087084",
  1178 => x"29bba005",
  1179 => x"7008e40c",
  1180 => x"5151bb98",
  1181 => x"08811187",
  1182 => x"06bb980c",
  1183 => x"51800bbb",
  1184 => x"cc0ca7bd",
  1185 => x"2da7c42d",
  1186 => x"0290050d",
  1187 => x"0402fc05",
  1188 => x"0da7ca2d",
  1189 => x"810bbbcc",
  1190 => x"0ca7c42d",
  1191 => x"bbcc0851",
  1192 => x"70fa3802",
  1193 => x"84050d04",
  1194 => x"02f8050d",
  1195 => x"baf051a1",
  1196 => x"c42da2d7",
  1197 => x"51a7b92d",
  1198 => x"a6e32d81",
  1199 => x"f452bb98",
  1200 => x"51a29b2d",
  1201 => x"0288050d",
  1202 => x"0402f405",
  1203 => x"0da6cb04",
  1204 => x"b5d00881",
  1205 => x"f02e0981",
  1206 => x"06893881",
  1207 => x"0bb5c40c",
  1208 => x"a6cb04b5",
  1209 => x"d00881e0",
  1210 => x"2e098106",
  1211 => x"8938810b",
  1212 => x"b5c80ca6",
  1213 => x"cb04b5d0",
  1214 => x"0852b5c8",
  1215 => x"08802e88",
  1216 => x"38b5d008",
  1217 => x"81800552",
  1218 => x"71842c72",
  1219 => x"8f065353",
  1220 => x"b5c40880",
  1221 => x"2e993872",
  1222 => x"8429b584",
  1223 => x"05721381",
  1224 => x"712b7009",
  1225 => x"73080673",
  1226 => x"0c515353",
  1227 => x"a6c10472",
  1228 => x"8429b584",
  1229 => x"05721383",
  1230 => x"712b7208",
  1231 => x"07720c53",
  1232 => x"53800bb5",
  1233 => x"c80c800b",
  1234 => x"b5c40cba",
  1235 => x"f051a1d7",
  1236 => x"2db5d008",
  1237 => x"ff24fef8",
  1238 => x"38800bb5",
  1239 => x"d00c028c",
  1240 => x"050d0402",
  1241 => x"f8050db5",
  1242 => x"84528f51",
  1243 => x"80727084",
  1244 => x"05540cff",
  1245 => x"11517080",
  1246 => x"25f23802",
  1247 => x"88050d04",
  1248 => x"02f0050d",
  1249 => x"7551a7ca",
  1250 => x"2d70822c",
  1251 => x"fc06b584",
  1252 => x"1172109e",
  1253 => x"06710870",
  1254 => x"722a7083",
  1255 => x"0682742b",
  1256 => x"70097406",
  1257 => x"760c5451",
  1258 => x"56575351",
  1259 => x"53a7c42d",
  1260 => x"71b5d00c",
  1261 => x"0290050d",
  1262 => x"0471980c",
  1263 => x"04ffb008",
  1264 => x"b5d00c04",
  1265 => x"810bffb0",
  1266 => x"0c04800b",
  1267 => x"ffb00c04",
  1268 => x"02fc050d",
  1269 => x"800bb5cc",
  1270 => x"0c805184",
  1271 => x"e52d0284",
  1272 => x"050d0402",
  1273 => x"f0050dbb",
  1274 => x"e4085481",
  1275 => x"f72d800b",
  1276 => x"bbe80c73",
  1277 => x"08802e80",
  1278 => x"eb38820b",
  1279 => x"b5e40cbb",
  1280 => x"e8088f06",
  1281 => x"b5e00c73",
  1282 => x"08527181",
  1283 => x"2ea43871",
  1284 => x"832e0981",
  1285 => x"06b93888",
  1286 => x"1480f52d",
  1287 => x"841508b3",
  1288 => x"84535452",
  1289 => x"85f32d71",
  1290 => x"84291370",
  1291 => x"085252a8",
  1292 => x"d304bbe0",
  1293 => x"08881508",
  1294 => x"2c708106",
  1295 => x"51527180",
  1296 => x"2e8738b3",
  1297 => x"8851a8cc",
  1298 => x"04b38c51",
  1299 => x"85f32d84",
  1300 => x"14085185",
  1301 => x"f32dbbe8",
  1302 => x"088105bb",
  1303 => x"e80c8c14",
  1304 => x"54a7f304",
  1305 => x"0290050d",
  1306 => x"0471bbe4",
  1307 => x"0ca7e32d",
  1308 => x"bbe808ff",
  1309 => x"05bbec0c",
  1310 => x"0402f005",
  1311 => x"0d8751a7",
  1312 => x"802db5d0",
  1313 => x"08812a70",
  1314 => x"81065152",
  1315 => x"71802ea0",
  1316 => x"38a99704",
  1317 => x"a5c92d87",
  1318 => x"51a7802d",
  1319 => x"b5d008f4",
  1320 => x"38b5cc08",
  1321 => x"813270b5",
  1322 => x"cc0c7052",
  1323 => x"5284e52d",
  1324 => x"b5cc0896",
  1325 => x"3880da51",
  1326 => x"a7802d81",
  1327 => x"f551a780",
  1328 => x"2d81f251",
  1329 => x"a7802dab",
  1330 => x"e70481f5",
  1331 => x"51a7802d",
  1332 => x"b5d00881",
  1333 => x"2a708106",
  1334 => x"51527180",
  1335 => x"2e8f38bb",
  1336 => x"ec085271",
  1337 => x"802e8638",
  1338 => x"ff12bbec",
  1339 => x"0c81f251",
  1340 => x"a7802db5",
  1341 => x"d008812a",
  1342 => x"70810651",
  1343 => x"5271802e",
  1344 => x"9538bbe8",
  1345 => x"08ff05bb",
  1346 => x"ec085452",
  1347 => x"72722586",
  1348 => x"388113bb",
  1349 => x"ec0c80da",
  1350 => x"51a7802d",
  1351 => x"b5d00881",
  1352 => x"2a708106",
  1353 => x"51527180",
  1354 => x"2e80fb38",
  1355 => x"bbe408bb",
  1356 => x"ec085553",
  1357 => x"73802e8a",
  1358 => x"388c13ff",
  1359 => x"155553aa",
  1360 => x"b4047208",
  1361 => x"5271822e",
  1362 => x"a6387182",
  1363 => x"26893871",
  1364 => x"812ea538",
  1365 => x"aba60471",
  1366 => x"832ead38",
  1367 => x"71842e09",
  1368 => x"810680c2",
  1369 => x"38881308",
  1370 => x"51a8e92d",
  1371 => x"aba60488",
  1372 => x"13085271",
  1373 => x"2daba604",
  1374 => x"810b8814",
  1375 => x"082bbbe0",
  1376 => x"0832bbe0",
  1377 => x"0caba304",
  1378 => x"881380f5",
  1379 => x"2d81058b",
  1380 => x"1480f52d",
  1381 => x"53547174",
  1382 => x"24833880",
  1383 => x"54738814",
  1384 => x"81b72da7",
  1385 => x"e32d8054",
  1386 => x"800bb5e4",
  1387 => x"0c738f06",
  1388 => x"b5e00ca0",
  1389 => x"5273bbec",
  1390 => x"082e0981",
  1391 => x"069838bb",
  1392 => x"e808ff05",
  1393 => x"74327009",
  1394 => x"81057072",
  1395 => x"079f2a91",
  1396 => x"71315151",
  1397 => x"53537151",
  1398 => x"82ee2d81",
  1399 => x"14548e74",
  1400 => x"25c638b5",
  1401 => x"cc085271",
  1402 => x"b5d00c02",
  1403 => x"90050d04",
  1404 => x"00ffffff",
  1405 => x"ff00ffff",
  1406 => x"ffff00ff",
  1407 => x"ffffff00",
  1408 => x"52657365",
  1409 => x"74000000",
  1410 => x"4f707469",
  1411 => x"6f6e7320",
  1412 => x"10000000",
  1413 => x"54757262",
  1414 => x"6f202831",
  1415 => x"302e3734",
  1416 => x"4d487a29",
  1417 => x"00000000",
  1418 => x"4d6f7573",
  1419 => x"6520656d",
  1420 => x"756c6174",
  1421 => x"696f6e00",
  1422 => x"45786974",
  1423 => x"00000000",
  1424 => x"5363616e",
  1425 => x"6c696e65",
  1426 => x"73000000",
  1427 => x"53442043",
  1428 => x"61726400",
  1429 => x"4a617061",
  1430 => x"6e657365",
  1431 => x"206b6579",
  1432 => x"626f6172",
  1433 => x"64206c61",
  1434 => x"796f7574",
  1435 => x"00000000",
  1436 => x"4261636b",
  1437 => x"00000000",
  1438 => x"32303438",
  1439 => x"4c422052",
  1440 => x"414d0000",
  1441 => x"34303936",
  1442 => x"4b422052",
  1443 => x"414d0000",
  1444 => x"536c323a",
  1445 => x"204e6f6e",
  1446 => x"65000000",
  1447 => x"536c323a",
  1448 => x"20455345",
  1449 => x"2d534343",
  1450 => x"20314d42",
  1451 => x"2f534343",
  1452 => x"2d490000",
  1453 => x"536c323a",
  1454 => x"20455345",
  1455 => x"2d52414d",
  1456 => x"20314d42",
  1457 => x"2f415343",
  1458 => x"49493800",
  1459 => x"536c323a",
  1460 => x"20455345",
  1461 => x"2d52414d",
  1462 => x"20314d42",
  1463 => x"2f415343",
  1464 => x"49493136",
  1465 => x"00000000",
  1466 => x"536c313a",
  1467 => x"204e6f6e",
  1468 => x"65000000",
  1469 => x"536c313a",
  1470 => x"20455345",
  1471 => x"2d534343",
  1472 => x"20314d42",
  1473 => x"2f534343",
  1474 => x"2d490000",
  1475 => x"536c313a",
  1476 => x"204d6567",
  1477 => x"6152414d",
  1478 => x"00000000",
  1479 => x"56474120",
  1480 => x"2d203331",
  1481 => x"4b487a2c",
  1482 => x"20363048",
  1483 => x"7a000000",
  1484 => x"56474120",
  1485 => x"2d203331",
  1486 => x"4b487a2c",
  1487 => x"20353048",
  1488 => x"7a000000",
  1489 => x"5456202d",
  1490 => x"20343830",
  1491 => x"692c2036",
  1492 => x"30487a00",
  1493 => x"496e6974",
  1494 => x"69616c69",
  1495 => x"7a696e67",
  1496 => x"20534420",
  1497 => x"63617264",
  1498 => x"0a000000",
  1499 => x"53444843",
  1500 => x"20636172",
  1501 => x"64206465",
  1502 => x"74656374",
  1503 => x"65642062",
  1504 => x"7574206e",
  1505 => x"6f740a73",
  1506 => x"7570706f",
  1507 => x"72746564",
  1508 => x"3b206469",
  1509 => x"7361626c",
  1510 => x"696e6720",
  1511 => x"53442063",
  1512 => x"6172640a",
  1513 => x"10204f4b",
  1514 => x"0a000000",
  1515 => x"46617433",
  1516 => x"32206669",
  1517 => x"6c657379",
  1518 => x"7374656d",
  1519 => x"20646574",
  1520 => x"65637465",
  1521 => x"64206275",
  1522 => x"740a6e6f",
  1523 => x"74207375",
  1524 => x"70706f72",
  1525 => x"7465643b",
  1526 => x"20646973",
  1527 => x"61626c69",
  1528 => x"6e672053",
  1529 => x"44206361",
  1530 => x"72640a10",
  1531 => x"204f4b0a",
  1532 => x"00000000",
  1533 => x"54727969",
  1534 => x"6e67204d",
  1535 => x"53583342",
  1536 => x"494f532e",
  1537 => x"5359532e",
  1538 => x"2e2e0a00",
  1539 => x"4d535833",
  1540 => x"42494f53",
  1541 => x"53595300",
  1542 => x"54727969",
  1543 => x"6e672042",
  1544 => x"494f535f",
  1545 => x"4d32502e",
  1546 => x"524f4d2e",
  1547 => x"2e2e0a00",
  1548 => x"42494f53",
  1549 => x"5f4d3250",
  1550 => x"524f4d00",
  1551 => x"4f70656e",
  1552 => x"65642042",
  1553 => x"494f532c",
  1554 => x"206c6f61",
  1555 => x"64696e67",
  1556 => x"2e2e2e0a",
  1557 => x"00000000",
  1558 => x"52656164",
  1559 => x"20626c6f",
  1560 => x"636b2066",
  1561 => x"61696c65",
  1562 => x"640a0000",
  1563 => x"4c6f6164",
  1564 => x"696e6720",
  1565 => x"42494f53",
  1566 => x"20666169",
  1567 => x"6c65640a",
  1568 => x"00000000",
  1569 => x"52656164",
  1570 => x"206f6620",
  1571 => x"4d425220",
  1572 => x"6661696c",
  1573 => x"65640a00",
  1574 => x"46415431",
  1575 => x"36202020",
  1576 => x"00000000",
  1577 => x"46415433",
  1578 => x"32202020",
  1579 => x"00000000",
  1580 => x"25642070",
  1581 => x"61727469",
  1582 => x"74696f6e",
  1583 => x"7320666f",
  1584 => x"756e640a",
  1585 => x"00000000",
  1586 => x"4e6f2070",
  1587 => x"61727469",
  1588 => x"74696f6e",
  1589 => x"20736967",
  1590 => x"6e617475",
  1591 => x"72652066",
  1592 => x"6f756e64",
  1593 => x"0a000000",
  1594 => x"556e7375",
  1595 => x"70706f72",
  1596 => x"74656420",
  1597 => x"70617274",
  1598 => x"6974696f",
  1599 => x"6e207479",
  1600 => x"7065210a",
  1601 => x"00000000",
  1602 => x"53444843",
  1603 => x"20496e69",
  1604 => x"7469616c",
  1605 => x"697a6174",
  1606 => x"696f6e20",
  1607 => x"6572726f",
  1608 => x"72210a00",
  1609 => x"434d4435",
  1610 => x"38202564",
  1611 => x"0a202000",
  1612 => x"496e6974",
  1613 => x"69616c69",
  1614 => x"7a696e67",
  1615 => x"20534420",
  1616 => x"63617264",
  1617 => x"2e2e2e0a",
  1618 => x"00000000",
  1619 => x"53442063",
  1620 => x"61726420",
  1621 => x"72657365",
  1622 => x"74206661",
  1623 => x"696c6564",
  1624 => x"210a0000",
  1625 => x"52656164",
  1626 => x"20636f6d",
  1627 => x"6d616e64",
  1628 => x"20666169",
  1629 => x"6c656420",
  1630 => x"61742025",
  1631 => x"64202825",
  1632 => x"64290a00",
  1633 => x"16200000",
  1634 => x"14200000",
  1635 => x"15200000",
  1636 => x"00000002",
  1637 => x"00000002",
  1638 => x"00001600",
  1639 => x"00000540",
  1640 => x"00000004",
  1641 => x"00001608",
  1642 => x"000019dc",
  1643 => x"00000001",
  1644 => x"00001614",
  1645 => x"00000007",
  1646 => x"00000001",
  1647 => x"00001628",
  1648 => x"0000000a",
  1649 => x"00000002",
  1650 => x"00001638",
  1651 => x"000013d0",
  1652 => x"00000000",
  1653 => x"00000000",
  1654 => x"00000000",
  1655 => x"00000003",
  1656 => x"00001a6c",
  1657 => x"00000003",
  1658 => x"00000001",
  1659 => x"00001640",
  1660 => x"0000000b",
  1661 => x"00000001",
  1662 => x"0000164c",
  1663 => x"00000002",
  1664 => x"00000003",
  1665 => x"00001a60",
  1666 => x"00000003",
  1667 => x"00000003",
  1668 => x"00001a50",
  1669 => x"00000004",
  1670 => x"00000001",
  1671 => x"00001654",
  1672 => x"00000006",
  1673 => x"00000003",
  1674 => x"00001a48",
  1675 => x"00000002",
  1676 => x"00000004",
  1677 => x"00001670",
  1678 => x"00001994",
  1679 => x"00000000",
  1680 => x"00000000",
  1681 => x"00000000",
  1682 => x"00001678",
  1683 => x"00001684",
  1684 => x"00001690",
  1685 => x"0000169c",
  1686 => x"000016b4",
  1687 => x"000016cc",
  1688 => x"000016e8",
  1689 => x"000016f4",
  1690 => x"0000170c",
  1691 => x"0000171c",
  1692 => x"00001730",
  1693 => x"00001744",
  1694 => x"00000003",
  1695 => x"00000000",
  1696 => x"00000000",
  1697 => x"00000000",
  1698 => x"00000000",
  1699 => x"00000000",
  1700 => x"00000000",
  1701 => x"00000000",
  1702 => x"00000000",
  1703 => x"00000000",
  1704 => x"00000000",
  1705 => x"00000000",
  1706 => x"00000000",
  1707 => x"00000000",
  1708 => x"00000000",
  1709 => x"00000000",
  1710 => x"00000000",
  1711 => x"00000000",
  1712 => x"00000000",
  1713 => x"00000000",
  1714 => x"00000000",
  1715 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

