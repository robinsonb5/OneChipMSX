-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b0bb4",
     9 => x"b0080b0b",
    10 => x"0bb4b408",
    11 => x"0b0b0bb4",
    12 => x"b8080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"b4b80c0b",
    16 => x"0b0bb4b4",
    17 => x"0c0b0b0b",
    18 => x"b4b00c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0baacc",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"b4b070ba",
    57 => x"90278b38",
    58 => x"80717084",
    59 => x"05530c81",
    60 => x"e2048c51",
    61 => x"8af10402",
    62 => x"fc050df8",
    63 => x"80518f0b",
    64 => x"b4c00c9f",
    65 => x"0bb4c40c",
    66 => x"a0717081",
    67 => x"055334b4",
    68 => x"c408ff05",
    69 => x"b4c40cb4",
    70 => x"c4088025",
    71 => x"eb38b4c0",
    72 => x"08ff05b4",
    73 => x"c00cb4c0",
    74 => x"088025d7",
    75 => x"38028405",
    76 => x"0d0402f0",
    77 => x"050df880",
    78 => x"53f8a054",
    79 => x"83bf5273",
    80 => x"70810555",
    81 => x"33517073",
    82 => x"70810555",
    83 => x"34ff1252",
    84 => x"718025eb",
    85 => x"38fbc053",
    86 => x"9f52a073",
    87 => x"70810555",
    88 => x"34ff1252",
    89 => x"718025f2",
    90 => x"38029005",
    91 => x"0d0402f4",
    92 => x"050d7453",
    93 => x"8e0bb4c0",
    94 => x"08258f38",
    95 => x"82b22db4",
    96 => x"c008ff05",
    97 => x"b4c00c82",
    98 => x"f404b4c0",
    99 => x"08b4c408",
   100 => x"5351728a",
   101 => x"2e098106",
   102 => x"b7387151",
   103 => x"719f24a0",
   104 => x"38b4c008",
   105 => x"a02911f8",
   106 => x"80115151",
   107 => x"a07134b4",
   108 => x"c4088105",
   109 => x"b4c40cb4",
   110 => x"c408519f",
   111 => x"7125e238",
   112 => x"800bb4c4",
   113 => x"0cb4c008",
   114 => x"8105b4c0",
   115 => x"0c83e404",
   116 => x"70a02912",
   117 => x"f8801151",
   118 => x"51727134",
   119 => x"b4c40881",
   120 => x"05b4c40c",
   121 => x"b4c408a0",
   122 => x"2e098106",
   123 => x"8e38800b",
   124 => x"b4c40cb4",
   125 => x"c0088105",
   126 => x"b4c00c02",
   127 => x"8c050d04",
   128 => x"02e8050d",
   129 => x"77795656",
   130 => x"880bfc16",
   131 => x"77712c8f",
   132 => x"06545254",
   133 => x"80537272",
   134 => x"25953871",
   135 => x"53fbe014",
   136 => x"51877134",
   137 => x"8114ff14",
   138 => x"545472f1",
   139 => x"387153f9",
   140 => x"1576712c",
   141 => x"87065351",
   142 => x"71802e8b",
   143 => x"38fbe014",
   144 => x"51717134",
   145 => x"81145472",
   146 => x"8e249538",
   147 => x"8f733153",
   148 => x"fbe01451",
   149 => x"a0713481",
   150 => x"14ff1454",
   151 => x"5472f138",
   152 => x"0298050d",
   153 => x"0402ec05",
   154 => x"0d800bb4",
   155 => x"c80cf68c",
   156 => x"08f69008",
   157 => x"71882c56",
   158 => x"5481ff06",
   159 => x"52737225",
   160 => x"88387154",
   161 => x"820bb4c8",
   162 => x"0c72882c",
   163 => x"7381ff06",
   164 => x"54557473",
   165 => x"258b3872",
   166 => x"b4c80884",
   167 => x"07b4c80c",
   168 => x"5573842b",
   169 => x"86a07125",
   170 => x"83713170",
   171 => x"0b0b0bb1",
   172 => x"9c0c8171",
   173 => x"2bff05f6",
   174 => x"880cfecc",
   175 => x"13ff122c",
   176 => x"788829ff",
   177 => x"94057081",
   178 => x"2cb4c808",
   179 => x"52585255",
   180 => x"51525476",
   181 => x"802e8538",
   182 => x"70810751",
   183 => x"70f6940c",
   184 => x"71098105",
   185 => x"f6800c72",
   186 => x"098105f6",
   187 => x"840c0294",
   188 => x"050d0402",
   189 => x"f4050d74",
   190 => x"53727081",
   191 => x"055480f5",
   192 => x"2d527180",
   193 => x"2e893871",
   194 => x"5182ee2d",
   195 => x"85f90402",
   196 => x"8c050d04",
   197 => x"02f8050d",
   198 => x"a2842d80",
   199 => x"da51a3bb",
   200 => x"2db4b008",
   201 => x"812a7081",
   202 => x"06515271",
   203 => x"802ee938",
   204 => x"0288050d",
   205 => x"0402f405",
   206 => x"0dba8008",
   207 => x"99c406b3",
   208 => x"8c0b80f5",
   209 => x"2d525270",
   210 => x"802e8638",
   211 => x"71848007",
   212 => x"52b2c40b",
   213 => x"80f52d72",
   214 => x"07b2dc0b",
   215 => x"80f52d70",
   216 => x"812a7081",
   217 => x"06515354",
   218 => x"5270802e",
   219 => x"86387182",
   220 => x"80075272",
   221 => x"81065170",
   222 => x"802e8538",
   223 => x"71880752",
   224 => x"b2e80b80",
   225 => x"f52d7084",
   226 => x"2b730781",
   227 => x"8432b4b0",
   228 => x"0c51028c",
   229 => x"050d0402",
   230 => x"f4050d74",
   231 => x"70818432",
   232 => x"ba800c70",
   233 => x"83065253",
   234 => x"70b2bc0b",
   235 => x"880581b7",
   236 => x"2d72892a",
   237 => x"70810651",
   238 => x"5170b38c",
   239 => x"0b81b72d",
   240 => x"72832a81",
   241 => x"0673882a",
   242 => x"70810651",
   243 => x"52527080",
   244 => x"2e853871",
   245 => x"82075271",
   246 => x"b2dc0b81",
   247 => x"b72d7284",
   248 => x"2c708306",
   249 => x"515170b2",
   250 => x"e80b81b7",
   251 => x"2d70b4b0",
   252 => x"0c028c05",
   253 => x"0d0402d4",
   254 => x"050dadd0",
   255 => x"5185f32d",
   256 => x"9af12db4",
   257 => x"b008802e",
   258 => x"82ab3886",
   259 => x"b52db4b0",
   260 => x"08538de0",
   261 => x"2db4b008",
   262 => x"54b4b008",
   263 => x"802e8297",
   264 => x"389dac2d",
   265 => x"b4b00880",
   266 => x"2e8738ad",
   267 => x"e85188be",
   268 => x"0496dd2d",
   269 => x"b4b00880",
   270 => x"2e9c38ae",
   271 => x"a85185f3",
   272 => x"2d86942d",
   273 => x"72840753",
   274 => x"810bfec4",
   275 => x"0c72fec0",
   276 => x"0c725187",
   277 => x"972d840b",
   278 => x"fec40cae",
   279 => x"f05185f3",
   280 => x"2daf8852",
   281 => x"b4d05193",
   282 => x"f22db4b0",
   283 => x"089838af",
   284 => x"945185f3",
   285 => x"2dafac52",
   286 => x"b4d05193",
   287 => x"f22db4b0",
   288 => x"08802e81",
   289 => x"b038afb8",
   290 => x"5185f32d",
   291 => x"b4d40857",
   292 => x"8077595a",
   293 => x"767a2e8b",
   294 => x"38811a78",
   295 => x"812a595a",
   296 => x"77f738f7",
   297 => x"1a5a8077",
   298 => x"25818038",
   299 => x"79527751",
   300 => x"84802db4",
   301 => x"dc52b4d0",
   302 => x"5196b72d",
   303 => x"b4b00853",
   304 => x"b4b00880",
   305 => x"2e80c938",
   306 => x"b4dc5b80",
   307 => x"5989fd04",
   308 => x"7a708405",
   309 => x"5c087081",
   310 => x"ff067188",
   311 => x"2c7081ff",
   312 => x"0673902c",
   313 => x"7081ff06",
   314 => x"75982afe",
   315 => x"c80cfec8",
   316 => x"0c58fec8",
   317 => x"0c57fec8",
   318 => x"0c841a5a",
   319 => x"53765384",
   320 => x"80772584",
   321 => x"38848053",
   322 => x"727924c4",
   323 => x"388a9b04",
   324 => x"afd45185",
   325 => x"f32d7254",
   326 => x"8ab704b4",
   327 => x"d051968a",
   328 => x"2dfc8017",
   329 => x"81195957",
   330 => x"89a60482",
   331 => x"0bfec40c",
   332 => x"81548ab7",
   333 => x"04805473",
   334 => x"b4b00c02",
   335 => x"ac050d04",
   336 => x"02f8050d",
   337 => x"a48b2d81",
   338 => x"f72d8151",
   339 => x"84e52dfe",
   340 => x"c4528172",
   341 => x"0ca1c82d",
   342 => x"a1c82d84",
   343 => x"720c87f6",
   344 => x"2db1a051",
   345 => x"a5e92d80",
   346 => x"5184e52d",
   347 => x"0288050d",
   348 => x"0402ec05",
   349 => x"0d8cb851",
   350 => x"87972d81",
   351 => x"0bfec40c",
   352 => x"8cb80bfe",
   353 => x"c00c840b",
   354 => x"fec40c83",
   355 => x"0bfecc0c",
   356 => x"a1e32da3",
   357 => x"ff2da1c8",
   358 => x"2da1c82d",
   359 => x"81f72d81",
   360 => x"5184e52d",
   361 => x"a1c82da1",
   362 => x"c82d8151",
   363 => x"84e52d87",
   364 => x"f62db4b0",
   365 => x"08802e81",
   366 => x"d4388051",
   367 => x"84e52db1",
   368 => x"a051a5e9",
   369 => x"2db9e808",
   370 => x"09708306",
   371 => x"fecc0c52",
   372 => x"b9e00889",
   373 => x"38b9e408",
   374 => x"802e80e2",
   375 => x"38fed008",
   376 => x"70810651",
   377 => x"5271802e",
   378 => x"80d438a4",
   379 => x"852db9e0",
   380 => x"0870b9e4",
   381 => x"08705755",
   382 => x"565280ff",
   383 => x"72258438",
   384 => x"80ff5280",
   385 => x"ff732584",
   386 => x"3880ff53",
   387 => x"71ff8025",
   388 => x"8438ff80",
   389 => x"5272ff80",
   390 => x"258438ff",
   391 => x"80537472",
   392 => x"31b9e00c",
   393 => x"737331b9",
   394 => x"e40ca3ff",
   395 => x"2d71882b",
   396 => x"83fe8006",
   397 => x"7381ff06",
   398 => x"7107fed0",
   399 => x"0c52a284",
   400 => x"2da5f92d",
   401 => x"b4b00853",
   402 => x"86b52db4",
   403 => x"b008fec0",
   404 => x"0c86b52d",
   405 => x"b4b008b4",
   406 => x"cc082e9c",
   407 => x"38b4b008",
   408 => x"b4cc0c84",
   409 => x"52725184",
   410 => x"e52da1c8",
   411 => x"2da1c82d",
   412 => x"ff125271",
   413 => x"8025ee38",
   414 => x"72802e89",
   415 => x"388a0bfe",
   416 => x"c40c8bc5",
   417 => x"04820bfe",
   418 => x"c40c8bc5",
   419 => x"04afe851",
   420 => x"85f32d82",
   421 => x"0bfec40c",
   422 => x"800bb4b0",
   423 => x"0c029405",
   424 => x"0d0402e8",
   425 => x"050d7779",
   426 => x"7b585555",
   427 => x"80537276",
   428 => x"25a33874",
   429 => x"70810556",
   430 => x"80f52d74",
   431 => x"70810556",
   432 => x"80f52d52",
   433 => x"5271712e",
   434 => x"86388151",
   435 => x"8dd70481",
   436 => x"13538dae",
   437 => x"04805170",
   438 => x"b4b00c02",
   439 => x"98050d04",
   440 => x"02d8050d",
   441 => x"800bb8e4",
   442 => x"0cb4dc52",
   443 => x"80519c91",
   444 => x"2db4b008",
   445 => x"54b4b008",
   446 => x"8c38b080",
   447 => x"5185f32d",
   448 => x"735592fb",
   449 => x"04805681",
   450 => x"0bb9880c",
   451 => x"8853b094",
   452 => x"52b59251",
   453 => x"8da22db4",
   454 => x"b008762e",
   455 => x"09810687",
   456 => x"38b4b008",
   457 => x"b9880c88",
   458 => x"53b0a052",
   459 => x"b5ae518d",
   460 => x"a22db4b0",
   461 => x"088738b4",
   462 => x"b008b988",
   463 => x"0cb98808",
   464 => x"802e80f6",
   465 => x"38b8a20b",
   466 => x"80f52db8",
   467 => x"a30b80f5",
   468 => x"2d71982b",
   469 => x"71902b07",
   470 => x"b8a40b80",
   471 => x"f52d7088",
   472 => x"2b7207b8",
   473 => x"a50b80f5",
   474 => x"2d7107b8",
   475 => x"da0b80f5",
   476 => x"2db8db0b",
   477 => x"80f52d71",
   478 => x"882b0753",
   479 => x"5f54525a",
   480 => x"56575573",
   481 => x"81abaa2e",
   482 => x"0981068d",
   483 => x"3875519d",
   484 => x"b32db4b0",
   485 => x"08568fa6",
   486 => x"047382d4",
   487 => x"d52e8738",
   488 => x"b0ac518f",
   489 => x"e704b4dc",
   490 => x"5275519c",
   491 => x"912db4b0",
   492 => x"0855b4b0",
   493 => x"08802e83",
   494 => x"c2388853",
   495 => x"b0a052b5",
   496 => x"ae518da2",
   497 => x"2db4b008",
   498 => x"8938810b",
   499 => x"b8e40c8f",
   500 => x"ed048853",
   501 => x"b09452b5",
   502 => x"92518da2",
   503 => x"2db4b008",
   504 => x"802e8a38",
   505 => x"b0c05185",
   506 => x"f32d90c7",
   507 => x"04b8da0b",
   508 => x"80f52d54",
   509 => x"7380d52e",
   510 => x"09810680",
   511 => x"ca38b8db",
   512 => x"0b80f52d",
   513 => x"547381aa",
   514 => x"2e098106",
   515 => x"ba38800b",
   516 => x"b4dc0b80",
   517 => x"f52d5654",
   518 => x"7481e92e",
   519 => x"83388154",
   520 => x"7481eb2e",
   521 => x"8c388055",
   522 => x"73752e09",
   523 => x"810682cb",
   524 => x"38b4e70b",
   525 => x"80f52d55",
   526 => x"748d38b4",
   527 => x"e80b80f5",
   528 => x"2d547382",
   529 => x"2e863880",
   530 => x"5592fb04",
   531 => x"b4e90b80",
   532 => x"f52d70b8",
   533 => x"dc0cff05",
   534 => x"b8e00cb4",
   535 => x"ea0b80f5",
   536 => x"2db4eb0b",
   537 => x"80f52d58",
   538 => x"76057782",
   539 => x"80290570",
   540 => x"b8e80cb4",
   541 => x"ec0b80f5",
   542 => x"2d70b8fc",
   543 => x"0cb8e408",
   544 => x"59575876",
   545 => x"802e81a3",
   546 => x"388853b0",
   547 => x"a052b5ae",
   548 => x"518da22d",
   549 => x"b4b00881",
   550 => x"e238b8dc",
   551 => x"0870842b",
   552 => x"b9800c70",
   553 => x"b8f80cb5",
   554 => x"810b80f5",
   555 => x"2db5800b",
   556 => x"80f52d71",
   557 => x"82802905",
   558 => x"b5820b80",
   559 => x"f52d7084",
   560 => x"80802912",
   561 => x"b5830b80",
   562 => x"f52d7081",
   563 => x"800a2912",
   564 => x"70b9840c",
   565 => x"b8fc0871",
   566 => x"29b8e808",
   567 => x"0570b8ec",
   568 => x"0cb5890b",
   569 => x"80f52db5",
   570 => x"880b80f5",
   571 => x"2d718280",
   572 => x"2905b58a",
   573 => x"0b80f52d",
   574 => x"70848080",
   575 => x"2912b58b",
   576 => x"0b80f52d",
   577 => x"70982b81",
   578 => x"f00a0672",
   579 => x"0570b8f0",
   580 => x"0cfe117e",
   581 => x"297705b8",
   582 => x"f40c5259",
   583 => x"5243545e",
   584 => x"51525952",
   585 => x"5d575957",
   586 => x"92f904b4",
   587 => x"ee0b80f5",
   588 => x"2db4ed0b",
   589 => x"80f52d71",
   590 => x"82802905",
   591 => x"70b9800c",
   592 => x"70a02983",
   593 => x"ff057089",
   594 => x"2a70b8f8",
   595 => x"0cb4f30b",
   596 => x"80f52db4",
   597 => x"f20b80f5",
   598 => x"2d718280",
   599 => x"290570b9",
   600 => x"840c7b71",
   601 => x"291e70b8",
   602 => x"f40c7db8",
   603 => x"f00c7305",
   604 => x"b8ec0c55",
   605 => x"5e515155",
   606 => x"55815574",
   607 => x"b4b00c02",
   608 => x"a8050d04",
   609 => x"02ec050d",
   610 => x"7670872c",
   611 => x"7180ff06",
   612 => x"555654b8",
   613 => x"e4088a38",
   614 => x"73882c74",
   615 => x"81ff0654",
   616 => x"55b4dc52",
   617 => x"b8e80815",
   618 => x"519c912d",
   619 => x"b4b00854",
   620 => x"b4b00880",
   621 => x"2eb338b8",
   622 => x"e408802e",
   623 => x"98387284",
   624 => x"29b4dc05",
   625 => x"70085253",
   626 => x"9db32db4",
   627 => x"b008f00a",
   628 => x"065393e7",
   629 => x"047210b4",
   630 => x"dc057080",
   631 => x"e02d5253",
   632 => x"9de32db4",
   633 => x"b0085372",
   634 => x"5473b4b0",
   635 => x"0c029405",
   636 => x"0d0402c8",
   637 => x"050d7f61",
   638 => x"5f5b800b",
   639 => x"b8f008b8",
   640 => x"f408595d",
   641 => x"56b8e408",
   642 => x"762e8a38",
   643 => x"b8dc0884",
   644 => x"2b58949b",
   645 => x"04b8f808",
   646 => x"842b5880",
   647 => x"59787827",
   648 => x"81a93878",
   649 => x"8f06a017",
   650 => x"5754738f",
   651 => x"38b4dc52",
   652 => x"76518117",
   653 => x"579c912d",
   654 => x"b4dc5680",
   655 => x"7680f52d",
   656 => x"56547474",
   657 => x"2e833881",
   658 => x"547481e5",
   659 => x"2e80f638",
   660 => x"81707506",
   661 => x"555d7380",
   662 => x"2e80ea38",
   663 => x"8b1680f5",
   664 => x"2d98065a",
   665 => x"7980de38",
   666 => x"8b537d52",
   667 => x"75518da2",
   668 => x"2db4b008",
   669 => x"80cf389c",
   670 => x"1608519d",
   671 => x"b32db4b0",
   672 => x"08841c0c",
   673 => x"9a1680e0",
   674 => x"2d519de3",
   675 => x"2db4b008",
   676 => x"b4b00888",
   677 => x"1d0cb4b0",
   678 => x"085555b8",
   679 => x"e408802e",
   680 => x"98389416",
   681 => x"80e02d51",
   682 => x"9de32db4",
   683 => x"b008902b",
   684 => x"83fff00a",
   685 => x"06701651",
   686 => x"5473881c",
   687 => x"0c797b0c",
   688 => x"7c549681",
   689 => x"04811959",
   690 => x"949d04b8",
   691 => x"e408802e",
   692 => x"ae387b51",
   693 => x"93842db4",
   694 => x"b008b4b0",
   695 => x"0880ffff",
   696 => x"fff80655",
   697 => x"5c7380ff",
   698 => x"fffff82e",
   699 => x"9238b4b0",
   700 => x"08fe05b8",
   701 => x"dc0829b8",
   702 => x"ec080557",
   703 => x"949b0480",
   704 => x"5473b4b0",
   705 => x"0c02b805",
   706 => x"0d0402f4",
   707 => x"050d7470",
   708 => x"08810571",
   709 => x"0c7008b8",
   710 => x"e0080653",
   711 => x"53718e38",
   712 => x"88130851",
   713 => x"93842db4",
   714 => x"b0088814",
   715 => x"0c810bb4",
   716 => x"b00c028c",
   717 => x"050d0402",
   718 => x"f0050d75",
   719 => x"881108fe",
   720 => x"05b8dc08",
   721 => x"29b8ec08",
   722 => x"117208b8",
   723 => x"e0080605",
   724 => x"79555354",
   725 => x"549c912d",
   726 => x"0290050d",
   727 => x"04b8e408",
   728 => x"b4b00c04",
   729 => x"02f4050d",
   730 => x"d45281ff",
   731 => x"720c7108",
   732 => x"5381ff72",
   733 => x"0c72882b",
   734 => x"83fe8006",
   735 => x"72087081",
   736 => x"ff065152",
   737 => x"5381ff72",
   738 => x"0c727107",
   739 => x"882b7208",
   740 => x"7081ff06",
   741 => x"51525381",
   742 => x"ff720c72",
   743 => x"7107882b",
   744 => x"72087081",
   745 => x"ff067207",
   746 => x"b4b00c52",
   747 => x"53028c05",
   748 => x"0d0402f4",
   749 => x"050d7476",
   750 => x"7181ff06",
   751 => x"d40c5353",
   752 => x"b98c0885",
   753 => x"3871892b",
   754 => x"5271982a",
   755 => x"d40c7190",
   756 => x"2a7081ff",
   757 => x"06d40c51",
   758 => x"71882a70",
   759 => x"81ff06d4",
   760 => x"0c517181",
   761 => x"ff06d40c",
   762 => x"72902a70",
   763 => x"81ff06d4",
   764 => x"0c51d408",
   765 => x"7081ff06",
   766 => x"515182b8",
   767 => x"bf527081",
   768 => x"ff2e0981",
   769 => x"06943881",
   770 => x"ff0bd40c",
   771 => x"d4087081",
   772 => x"ff06ff14",
   773 => x"54515171",
   774 => x"e53870b4",
   775 => x"b00c028c",
   776 => x"050d0402",
   777 => x"fc050d81",
   778 => x"c75181ff",
   779 => x"0bd40cff",
   780 => x"11517080",
   781 => x"25f43802",
   782 => x"84050d04",
   783 => x"02f0050d",
   784 => x"98a32d8f",
   785 => x"cf538052",
   786 => x"87fc80f7",
   787 => x"5197b22d",
   788 => x"b4b00854",
   789 => x"b4b00881",
   790 => x"2e098106",
   791 => x"a33881ff",
   792 => x"0bd40c82",
   793 => x"0a52849c",
   794 => x"80e95197",
   795 => x"b22db4b0",
   796 => x"088b3881",
   797 => x"ff0bd40c",
   798 => x"73539986",
   799 => x"0498a32d",
   800 => x"ff135372",
   801 => x"c13872b4",
   802 => x"b00c0290",
   803 => x"050d0402",
   804 => x"f4050d81",
   805 => x"ff0bd40c",
   806 => x"93538052",
   807 => x"87fc80c1",
   808 => x"5197b22d",
   809 => x"b4b0088b",
   810 => x"3881ff0b",
   811 => x"d40c8153",
   812 => x"99bc0498",
   813 => x"a32dff13",
   814 => x"5372df38",
   815 => x"72b4b00c",
   816 => x"028c050d",
   817 => x"0402f005",
   818 => x"0d98a32d",
   819 => x"83aa5284",
   820 => x"9c80c851",
   821 => x"97b22db4",
   822 => x"b008812e",
   823 => x"09810692",
   824 => x"3896e42d",
   825 => x"b4b00883",
   826 => x"ffff0653",
   827 => x"7283aa2e",
   828 => x"9738998f",
   829 => x"2d9a8304",
   830 => x"81549ae8",
   831 => x"04b0cc51",
   832 => x"85f32d80",
   833 => x"549ae804",
   834 => x"81ff0bd4",
   835 => x"0cb15398",
   836 => x"bc2db4b0",
   837 => x"08802e80",
   838 => x"c0388052",
   839 => x"87fc80fa",
   840 => x"5197b22d",
   841 => x"b4b008b1",
   842 => x"3881ff0b",
   843 => x"d40cd408",
   844 => x"5381ff0b",
   845 => x"d40c81ff",
   846 => x"0bd40c81",
   847 => x"ff0bd40c",
   848 => x"81ff0bd4",
   849 => x"0c72862a",
   850 => x"708106b4",
   851 => x"b0085651",
   852 => x"5372802e",
   853 => x"933899f8",
   854 => x"0472822e",
   855 => x"ff9f38ff",
   856 => x"135372ff",
   857 => x"aa387254",
   858 => x"73b4b00c",
   859 => x"0290050d",
   860 => x"0402f405",
   861 => x"0d810bb9",
   862 => x"8c0cd008",
   863 => x"708f2a70",
   864 => x"81065151",
   865 => x"5372f338",
   866 => x"72d00c98",
   867 => x"a32db0dc",
   868 => x"5185f32d",
   869 => x"d008708f",
   870 => x"2a708106",
   871 => x"51515372",
   872 => x"f338810b",
   873 => x"d00c80e3",
   874 => x"53805284",
   875 => x"d480c051",
   876 => x"97b22db4",
   877 => x"b008812e",
   878 => x"9a387282",
   879 => x"2e098106",
   880 => x"8c38b0e8",
   881 => x"5185f32d",
   882 => x"80539c88",
   883 => x"04ff1353",
   884 => x"72d73899",
   885 => x"c52db4b0",
   886 => x"08b98c0c",
   887 => x"b4b0088b",
   888 => x"38815287",
   889 => x"fc80d051",
   890 => x"97b22d81",
   891 => x"ff0bd40c",
   892 => x"d008708f",
   893 => x"2a708106",
   894 => x"51515372",
   895 => x"f33872d0",
   896 => x"0c81ff0b",
   897 => x"d40c8153",
   898 => x"72b4b00c",
   899 => x"028c050d",
   900 => x"0402e805",
   901 => x"0d785580",
   902 => x"5681ff0b",
   903 => x"d40cd008",
   904 => x"708f2a70",
   905 => x"81065151",
   906 => x"5372f338",
   907 => x"82810bd0",
   908 => x"0c81ff0b",
   909 => x"d40c7752",
   910 => x"87fc80d1",
   911 => x"5197b22d",
   912 => x"80dbc6df",
   913 => x"54b4b008",
   914 => x"802e8a38",
   915 => x"b1805185",
   916 => x"f32d9da3",
   917 => x"0481ff0b",
   918 => x"d40cd408",
   919 => x"7081ff06",
   920 => x"51537281",
   921 => x"fe2e0981",
   922 => x"069d3880",
   923 => x"ff5396e4",
   924 => x"2db4b008",
   925 => x"75708405",
   926 => x"570cff13",
   927 => x"53728025",
   928 => x"ed388156",
   929 => x"9d8d04ff",
   930 => x"145473c9",
   931 => x"3881ff0b",
   932 => x"d40cd008",
   933 => x"708f2a70",
   934 => x"81065151",
   935 => x"5372f338",
   936 => x"72d00c75",
   937 => x"b4b00c02",
   938 => x"98050d04",
   939 => x"b98c08b4",
   940 => x"b00c0402",
   941 => x"f4050d74",
   942 => x"70882a83",
   943 => x"fe800670",
   944 => x"72982a07",
   945 => x"72882b87",
   946 => x"fc808006",
   947 => x"73982b81",
   948 => x"f00a0671",
   949 => x"730707b4",
   950 => x"b00c5651",
   951 => x"5351028c",
   952 => x"050d0402",
   953 => x"f8050d02",
   954 => x"8e0580f5",
   955 => x"2d74882b",
   956 => x"077083ff",
   957 => x"ff06b4b0",
   958 => x"0c510288",
   959 => x"050d0402",
   960 => x"fc050d72",
   961 => x"5180710c",
   962 => x"800b8412",
   963 => x"0c028405",
   964 => x"0d0402f0",
   965 => x"050d7570",
   966 => x"08841208",
   967 => x"535353ff",
   968 => x"5471712e",
   969 => x"a838a485",
   970 => x"2d841308",
   971 => x"70842914",
   972 => x"88117008",
   973 => x"7081ff06",
   974 => x"84180881",
   975 => x"11870684",
   976 => x"1a0c5351",
   977 => x"55515151",
   978 => x"a3ff2d71",
   979 => x"5473b4b0",
   980 => x"0c029005",
   981 => x"0d0402f4",
   982 => x"050d7453",
   983 => x"84130881",
   984 => x"11870674",
   985 => x"08545151",
   986 => x"71712ef0",
   987 => x"38a4852d",
   988 => x"84130870",
   989 => x"84291488",
   990 => x"1178710c",
   991 => x"51515184",
   992 => x"13088111",
   993 => x"87068415",
   994 => x"0c51a3ff",
   995 => x"2d028c05",
   996 => x"0d0402f0",
   997 => x"050da485",
   998 => x"2de008e4",
   999 => x"08718b2a",
  1000 => x"70810651",
  1001 => x"53555270",
  1002 => x"802e9d38",
  1003 => x"b9900870",
  1004 => x"8429b998",
  1005 => x"057381ff",
  1006 => x"06710c51",
  1007 => x"51b99008",
  1008 => x"81118706",
  1009 => x"b9900c51",
  1010 => x"738b2a70",
  1011 => x"81065151",
  1012 => x"70802e81",
  1013 => x"8938b3e0",
  1014 => x"088429b9",
  1015 => x"f0057481",
  1016 => x"ff06710c",
  1017 => x"51b3e008",
  1018 => x"8105b3e0",
  1019 => x"0c850bb3",
  1020 => x"dc0cb3e0",
  1021 => x"08b3d808",
  1022 => x"2e098106",
  1023 => x"81863880",
  1024 => x"0bb3e00c",
  1025 => x"b9f00870",
  1026 => x"8306b9e8",
  1027 => x"0c70852a",
  1028 => x"708106b9",
  1029 => x"e4085651",
  1030 => x"52527080",
  1031 => x"2e8e38b9",
  1032 => x"f808fe80",
  1033 => x"3213b9e4",
  1034 => x"0ca0b304",
  1035 => x"b9f80813",
  1036 => x"b9e40c71",
  1037 => x"842a7081",
  1038 => x"06b9e008",
  1039 => x"54515170",
  1040 => x"802e9038",
  1041 => x"b9f40881",
  1042 => x"ff321281",
  1043 => x"05b9e00c",
  1044 => x"a1840471",
  1045 => x"b9f40831",
  1046 => x"b9e00ca1",
  1047 => x"8404b3dc",
  1048 => x"08ff05b3",
  1049 => x"dc0cb3dc",
  1050 => x"08ff2e09",
  1051 => x"81069538",
  1052 => x"b3e00880",
  1053 => x"2e8a3887",
  1054 => x"0bb3d808",
  1055 => x"31b3d80c",
  1056 => x"70b3e00c",
  1057 => x"738a2a70",
  1058 => x"81065151",
  1059 => x"70802ea8",
  1060 => x"38b9b808",
  1061 => x"b9bc0852",
  1062 => x"5271712e",
  1063 => x"9b38b9b8",
  1064 => x"08708429",
  1065 => x"b9c00570",
  1066 => x"08e40c51",
  1067 => x"51b9b808",
  1068 => x"81118706",
  1069 => x"b9b80c51",
  1070 => x"800bb9ec",
  1071 => x"0ca3f82d",
  1072 => x"a3ff2d02",
  1073 => x"90050d04",
  1074 => x"02fc050d",
  1075 => x"a4852d81",
  1076 => x"0bb9ec0c",
  1077 => x"a3ff2db9",
  1078 => x"ec085170",
  1079 => x"fa380284",
  1080 => x"050d0402",
  1081 => x"f8050db9",
  1082 => x"90519dff",
  1083 => x"2d9f9251",
  1084 => x"a3f42da3",
  1085 => x"9e2d81f4",
  1086 => x"52b9b851",
  1087 => x"9ed62d02",
  1088 => x"88050d04",
  1089 => x"02f4050d",
  1090 => x"a38604b4",
  1091 => x"b00881f0",
  1092 => x"2e098106",
  1093 => x"8938810b",
  1094 => x"b4a40ca3",
  1095 => x"8604b4b0",
  1096 => x"0881e02e",
  1097 => x"09810689",
  1098 => x"38810bb4",
  1099 => x"a80ca386",
  1100 => x"04b4b008",
  1101 => x"52b4a808",
  1102 => x"802e8838",
  1103 => x"b4b00881",
  1104 => x"80055271",
  1105 => x"842c728f",
  1106 => x"065353b4",
  1107 => x"a408802e",
  1108 => x"99387284",
  1109 => x"29b3e405",
  1110 => x"72138171",
  1111 => x"2b700973",
  1112 => x"0806730c",
  1113 => x"515353a2",
  1114 => x"fc047284",
  1115 => x"29b3e405",
  1116 => x"72138371",
  1117 => x"2b720807",
  1118 => x"720c5353",
  1119 => x"800bb4a8",
  1120 => x"0c800bb4",
  1121 => x"a40cb990",
  1122 => x"519e922d",
  1123 => x"b4b008ff",
  1124 => x"24fef838",
  1125 => x"800bb4b0",
  1126 => x"0c028c05",
  1127 => x"0d0402f8",
  1128 => x"050db3e4",
  1129 => x"528f5180",
  1130 => x"72708405",
  1131 => x"540cff11",
  1132 => x"51708025",
  1133 => x"f2380288",
  1134 => x"050d0402",
  1135 => x"f0050d75",
  1136 => x"51a4852d",
  1137 => x"70822cfc",
  1138 => x"06b3e411",
  1139 => x"72109e06",
  1140 => x"71087072",
  1141 => x"2a708306",
  1142 => x"82742b70",
  1143 => x"09740676",
  1144 => x"0c545156",
  1145 => x"57535153",
  1146 => x"a3ff2d71",
  1147 => x"b4b00c02",
  1148 => x"90050d04",
  1149 => x"71980c04",
  1150 => x"ffb008b4",
  1151 => x"b00c0481",
  1152 => x"0bffb00c",
  1153 => x"04800bff",
  1154 => x"b00c0402",
  1155 => x"fc050d80",
  1156 => x"0bb4ac0c",
  1157 => x"805184e5",
  1158 => x"2d028405",
  1159 => x"0d0402ec",
  1160 => x"050d7654",
  1161 => x"8052870b",
  1162 => x"881580f5",
  1163 => x"2d565374",
  1164 => x"72248338",
  1165 => x"a0537251",
  1166 => x"82ee2d81",
  1167 => x"128b1580",
  1168 => x"f52d5452",
  1169 => x"727225de",
  1170 => x"38029405",
  1171 => x"0d0402f0",
  1172 => x"050dba84",
  1173 => x"085481f7",
  1174 => x"2d800bba",
  1175 => x"880c7308",
  1176 => x"802e8180",
  1177 => x"38820bb4",
  1178 => x"c40cba88",
  1179 => x"088f06b4",
  1180 => x"c00c7308",
  1181 => x"5271832e",
  1182 => x"96387183",
  1183 => x"26893871",
  1184 => x"812eaf38",
  1185 => x"a5cf0471",
  1186 => x"852e9f38",
  1187 => x"a5cf0488",
  1188 => x"1480f52d",
  1189 => x"841508b1",
  1190 => x"90535452",
  1191 => x"85f32d71",
  1192 => x"84291370",
  1193 => x"085252a5",
  1194 => x"d3047351",
  1195 => x"a49e2da5",
  1196 => x"cf04ba80",
  1197 => x"08881508",
  1198 => x"2c708106",
  1199 => x"51527180",
  1200 => x"2e8738b1",
  1201 => x"9451a5cc",
  1202 => x"04b19851",
  1203 => x"85f32d84",
  1204 => x"14085185",
  1205 => x"f32dba88",
  1206 => x"088105ba",
  1207 => x"880c8c14",
  1208 => x"54a4de04",
  1209 => x"0290050d",
  1210 => x"0471ba84",
  1211 => x"0ca4ce2d",
  1212 => x"ba8808ff",
  1213 => x"05ba8c0c",
  1214 => x"0402ec05",
  1215 => x"0dba8408",
  1216 => x"5580f851",
  1217 => x"a3bb2db4",
  1218 => x"b008812a",
  1219 => x"70810651",
  1220 => x"52719b38",
  1221 => x"8751a3bb",
  1222 => x"2db4b008",
  1223 => x"812a7081",
  1224 => x"06515271",
  1225 => x"802eb138",
  1226 => x"a6ae04a2",
  1227 => x"842d8751",
  1228 => x"a3bb2db4",
  1229 => x"b008f438",
  1230 => x"a6be04a2",
  1231 => x"842d80f8",
  1232 => x"51a3bb2d",
  1233 => x"b4b008f3",
  1234 => x"38b4ac08",
  1235 => x"813270b4",
  1236 => x"ac0c7052",
  1237 => x"5284e52d",
  1238 => x"b4ac08a2",
  1239 => x"3880da51",
  1240 => x"a3bb2d81",
  1241 => x"f551a3bb",
  1242 => x"2d81f251",
  1243 => x"a3bb2d81",
  1244 => x"eb51a3bb",
  1245 => x"2d81f451",
  1246 => x"a3bb2daa",
  1247 => x"c20481f5",
  1248 => x"51a3bb2d",
  1249 => x"b4b00881",
  1250 => x"2a708106",
  1251 => x"51527180",
  1252 => x"2e8f38ba",
  1253 => x"8c085271",
  1254 => x"802e8638",
  1255 => x"ff12ba8c",
  1256 => x"0c81f251",
  1257 => x"a3bb2db4",
  1258 => x"b008812a",
  1259 => x"70810651",
  1260 => x"5271802e",
  1261 => x"9538ba88",
  1262 => x"08ff05ba",
  1263 => x"8c085452",
  1264 => x"72722586",
  1265 => x"388113ba",
  1266 => x"8c0cba8c",
  1267 => x"08705354",
  1268 => x"73802e8a",
  1269 => x"388c15ff",
  1270 => x"155555a7",
  1271 => x"d004820b",
  1272 => x"b4c40c71",
  1273 => x"8f06b4c0",
  1274 => x"0c81eb51",
  1275 => x"a3bb2db4",
  1276 => x"b008812a",
  1277 => x"70810651",
  1278 => x"5271802e",
  1279 => x"ad387408",
  1280 => x"852e0981",
  1281 => x"06a43888",
  1282 => x"1580f52d",
  1283 => x"ff055271",
  1284 => x"881681b7",
  1285 => x"2d71982b",
  1286 => x"52718025",
  1287 => x"8838800b",
  1288 => x"881681b7",
  1289 => x"2d7451a4",
  1290 => x"9e2d81f4",
  1291 => x"51a3bb2d",
  1292 => x"b4b00881",
  1293 => x"2a708106",
  1294 => x"51527180",
  1295 => x"2eb33874",
  1296 => x"08852e09",
  1297 => x"8106aa38",
  1298 => x"881580f5",
  1299 => x"2d810552",
  1300 => x"71881681",
  1301 => x"b72d7181",
  1302 => x"ff068b16",
  1303 => x"80f52d54",
  1304 => x"52727227",
  1305 => x"87387288",
  1306 => x"1681b72d",
  1307 => x"7451a49e",
  1308 => x"2d80da51",
  1309 => x"a3bb2db4",
  1310 => x"b008812a",
  1311 => x"70810651",
  1312 => x"5271802e",
  1313 => x"80fb38ba",
  1314 => x"8408ba8c",
  1315 => x"08555373",
  1316 => x"802e8a38",
  1317 => x"8c13ff15",
  1318 => x"5553a98f",
  1319 => x"04720852",
  1320 => x"71822ea6",
  1321 => x"38718226",
  1322 => x"89387181",
  1323 => x"2ea538aa",
  1324 => x"81047183",
  1325 => x"2ead3871",
  1326 => x"842e0981",
  1327 => x"0680c238",
  1328 => x"88130851",
  1329 => x"a5e92daa",
  1330 => x"81048813",
  1331 => x"0852712d",
  1332 => x"aa810481",
  1333 => x"0b881408",
  1334 => x"2bba8008",
  1335 => x"32ba800c",
  1336 => x"a9fe0488",
  1337 => x"1380f52d",
  1338 => x"81058b14",
  1339 => x"80f52d53",
  1340 => x"54717424",
  1341 => x"83388054",
  1342 => x"73881481",
  1343 => x"b72da4ce",
  1344 => x"2d805480",
  1345 => x"0bb4c40c",
  1346 => x"738f06b4",
  1347 => x"c00ca052",
  1348 => x"73ba8c08",
  1349 => x"2e098106",
  1350 => x"9838ba88",
  1351 => x"08ff0574",
  1352 => x"32700981",
  1353 => x"05707207",
  1354 => x"9f2a9171",
  1355 => x"31515153",
  1356 => x"53715182",
  1357 => x"ee2d8114",
  1358 => x"548e7425",
  1359 => x"c638b4ac",
  1360 => x"085271b4",
  1361 => x"b00c0294",
  1362 => x"050d0400",
  1363 => x"00ffffff",
  1364 => x"ff00ffff",
  1365 => x"ffff00ff",
  1366 => x"ffffff00",
  1367 => x"52657365",
  1368 => x"74000000",
  1369 => x"4f707469",
  1370 => x"6f6e7320",
  1371 => x"10000000",
  1372 => x"536f756e",
  1373 => x"64201000",
  1374 => x"54757262",
  1375 => x"6f202831",
  1376 => x"302e3734",
  1377 => x"4d487a29",
  1378 => x"00000000",
  1379 => x"4d6f7573",
  1380 => x"6520656d",
  1381 => x"756c6174",
  1382 => x"696f6e00",
  1383 => x"45786974",
  1384 => x"00000000",
  1385 => x"4d617374",
  1386 => x"65720000",
  1387 => x"4f504c4c",
  1388 => x"00000000",
  1389 => x"53434300",
  1390 => x"50534700",
  1391 => x"4261636b",
  1392 => x"00000000",
  1393 => x"5363616e",
  1394 => x"6c696e65",
  1395 => x"73000000",
  1396 => x"53442043",
  1397 => x"61726400",
  1398 => x"4a617061",
  1399 => x"6e657365",
  1400 => x"206b6579",
  1401 => x"626f6172",
  1402 => x"64206c61",
  1403 => x"796f7574",
  1404 => x"00000000",
  1405 => x"32303438",
  1406 => x"4c422052",
  1407 => x"414d0000",
  1408 => x"34303936",
  1409 => x"4b422052",
  1410 => x"414d0000",
  1411 => x"536c323a",
  1412 => x"204e6f6e",
  1413 => x"65000000",
  1414 => x"536c323a",
  1415 => x"20455345",
  1416 => x"2d534343",
  1417 => x"20314d42",
  1418 => x"2f534343",
  1419 => x"2d490000",
  1420 => x"536c323a",
  1421 => x"20455345",
  1422 => x"2d52414d",
  1423 => x"20314d42",
  1424 => x"2f415343",
  1425 => x"49493800",
  1426 => x"536c323a",
  1427 => x"20455345",
  1428 => x"2d52414d",
  1429 => x"20314d42",
  1430 => x"2f415343",
  1431 => x"49493136",
  1432 => x"00000000",
  1433 => x"536c313a",
  1434 => x"204e6f6e",
  1435 => x"65000000",
  1436 => x"536c313a",
  1437 => x"20455345",
  1438 => x"2d534343",
  1439 => x"20314d42",
  1440 => x"2f534343",
  1441 => x"2d490000",
  1442 => x"536c313a",
  1443 => x"204d6567",
  1444 => x"6152414d",
  1445 => x"00000000",
  1446 => x"56474120",
  1447 => x"2d203331",
  1448 => x"4b487a2c",
  1449 => x"20363048",
  1450 => x"7a000000",
  1451 => x"56474120",
  1452 => x"2d203331",
  1453 => x"4b487a2c",
  1454 => x"20353048",
  1455 => x"7a000000",
  1456 => x"5456202d",
  1457 => x"20343830",
  1458 => x"692c2036",
  1459 => x"30487a00",
  1460 => x"496e6974",
  1461 => x"69616c69",
  1462 => x"7a696e67",
  1463 => x"20534420",
  1464 => x"63617264",
  1465 => x"0a000000",
  1466 => x"53444843",
  1467 => x"20636172",
  1468 => x"64206465",
  1469 => x"74656374",
  1470 => x"65642062",
  1471 => x"7574206e",
  1472 => x"6f740a73",
  1473 => x"7570706f",
  1474 => x"72746564",
  1475 => x"3b206469",
  1476 => x"7361626c",
  1477 => x"696e6720",
  1478 => x"53442063",
  1479 => x"6172640a",
  1480 => x"10204f4b",
  1481 => x"0a000000",
  1482 => x"46617433",
  1483 => x"32206669",
  1484 => x"6c657379",
  1485 => x"7374656d",
  1486 => x"20646574",
  1487 => x"65637465",
  1488 => x"64206275",
  1489 => x"740a6e6f",
  1490 => x"74207375",
  1491 => x"70706f72",
  1492 => x"7465643b",
  1493 => x"20646973",
  1494 => x"61626c69",
  1495 => x"6e672053",
  1496 => x"44206361",
  1497 => x"72640a10",
  1498 => x"204f4b0a",
  1499 => x"00000000",
  1500 => x"54727969",
  1501 => x"6e67204d",
  1502 => x"53583342",
  1503 => x"494f532e",
  1504 => x"5359532e",
  1505 => x"2e2e0a00",
  1506 => x"4d535833",
  1507 => x"42494f53",
  1508 => x"53595300",
  1509 => x"54727969",
  1510 => x"6e672042",
  1511 => x"494f535f",
  1512 => x"4d32502e",
  1513 => x"524f4d2e",
  1514 => x"2e2e0a00",
  1515 => x"42494f53",
  1516 => x"5f4d3250",
  1517 => x"524f4d00",
  1518 => x"4f70656e",
  1519 => x"65642042",
  1520 => x"494f532c",
  1521 => x"206c6f61",
  1522 => x"64696e67",
  1523 => x"2e2e2e0a",
  1524 => x"00000000",
  1525 => x"52656164",
  1526 => x"20626c6f",
  1527 => x"636b2066",
  1528 => x"61696c65",
  1529 => x"640a0000",
  1530 => x"4c6f6164",
  1531 => x"696e6720",
  1532 => x"42494f53",
  1533 => x"20666169",
  1534 => x"6c65640a",
  1535 => x"00000000",
  1536 => x"52656164",
  1537 => x"206f6620",
  1538 => x"4d425220",
  1539 => x"6661696c",
  1540 => x"65640a00",
  1541 => x"46415431",
  1542 => x"36202020",
  1543 => x"00000000",
  1544 => x"46415433",
  1545 => x"32202020",
  1546 => x"00000000",
  1547 => x"4e6f2070",
  1548 => x"61727469",
  1549 => x"74696f6e",
  1550 => x"20736967",
  1551 => x"0a000000",
  1552 => x"42616420",
  1553 => x"70617274",
  1554 => x"0a000000",
  1555 => x"53444843",
  1556 => x"20657272",
  1557 => x"6f72210a",
  1558 => x"00000000",
  1559 => x"53442069",
  1560 => x"6e69742e",
  1561 => x"2e2e0a00",
  1562 => x"53442063",
  1563 => x"61726420",
  1564 => x"72657365",
  1565 => x"74206661",
  1566 => x"696c6564",
  1567 => x"210a0000",
  1568 => x"52656164",
  1569 => x"20666169",
  1570 => x"6c65640a",
  1571 => x"00000000",
  1572 => x"16200000",
  1573 => x"14200000",
  1574 => x"15200000",
  1575 => x"00000002",
  1576 => x"00000002",
  1577 => x"0000155c",
  1578 => x"00000540",
  1579 => x"00000004",
  1580 => x"00001564",
  1581 => x"0000193c",
  1582 => x"00000004",
  1583 => x"00001570",
  1584 => x"000018f4",
  1585 => x"00000001",
  1586 => x"00001578",
  1587 => x"00000007",
  1588 => x"00000001",
  1589 => x"0000158c",
  1590 => x"0000000a",
  1591 => x"00000002",
  1592 => x"0000159c",
  1593 => x"0000120b",
  1594 => x"00000000",
  1595 => x"00000000",
  1596 => x"00000000",
  1597 => x"00000005",
  1598 => x"000015a4",
  1599 => x"00000007",
  1600 => x"00000005",
  1601 => x"000015ac",
  1602 => x"00000007",
  1603 => x"00000005",
  1604 => x"000015b4",
  1605 => x"00000007",
  1606 => x"00000005",
  1607 => x"000015b8",
  1608 => x"00000007",
  1609 => x"00000004",
  1610 => x"000015bc",
  1611 => x"000018a0",
  1612 => x"00000000",
  1613 => x"00000000",
  1614 => x"00000000",
  1615 => x"00000003",
  1616 => x"000019cc",
  1617 => x"00000003",
  1618 => x"00000001",
  1619 => x"000015c4",
  1620 => x"0000000b",
  1621 => x"00000001",
  1622 => x"000015d0",
  1623 => x"00000002",
  1624 => x"00000003",
  1625 => x"000019c0",
  1626 => x"00000003",
  1627 => x"00000003",
  1628 => x"000019b0",
  1629 => x"00000004",
  1630 => x"00000001",
  1631 => x"000015d8",
  1632 => x"00000006",
  1633 => x"00000003",
  1634 => x"000019a8",
  1635 => x"00000002",
  1636 => x"00000004",
  1637 => x"000015bc",
  1638 => x"000018a0",
  1639 => x"00000000",
  1640 => x"00000000",
  1641 => x"00000000",
  1642 => x"000015f4",
  1643 => x"00001600",
  1644 => x"0000160c",
  1645 => x"00001618",
  1646 => x"00001630",
  1647 => x"00001648",
  1648 => x"00001664",
  1649 => x"00001670",
  1650 => x"00001688",
  1651 => x"00001698",
  1652 => x"000016ac",
  1653 => x"000016c0",
  1654 => x"00000003",
  1655 => x"00000000",
  1656 => x"00000000",
  1657 => x"00000000",
  1658 => x"00000000",
  1659 => x"00000000",
  1660 => x"00000000",
  1661 => x"00000000",
  1662 => x"00000000",
  1663 => x"00000000",
  1664 => x"00000000",
  1665 => x"00000000",
  1666 => x"00000000",
  1667 => x"00000000",
  1668 => x"00000000",
  1669 => x"00000000",
  1670 => x"00000000",
  1671 => x"00000000",
  1672 => x"00000000",
  1673 => x"00000000",
  1674 => x"00000000",
  1675 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

