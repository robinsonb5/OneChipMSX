-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b0bb0",
     9 => x"c4080b0b",
    10 => x"0bb0c808",
    11 => x"0b0b0bb0",
    12 => x"cc080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"b0cc0c0b",
    16 => x"0b0bb0c8",
    17 => x"0c0b0b0b",
    18 => x"b0c40c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0ba794",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"b0c470b6",
    57 => x"a0278b38",
    58 => x"80717084",
    59 => x"05530c81",
    60 => x"e2048c51",
    61 => x"87f20402",
    62 => x"fc050df8",
    63 => x"80518f0b",
    64 => x"b0d40c9f",
    65 => x"0bb0d80c",
    66 => x"a0717081",
    67 => x"055334b0",
    68 => x"d808ff05",
    69 => x"b0d80cb0",
    70 => x"d8088025",
    71 => x"eb38b0d4",
    72 => x"08ff05b0",
    73 => x"d40cb0d4",
    74 => x"088025d7",
    75 => x"38028405",
    76 => x"0d0402f0",
    77 => x"050df880",
    78 => x"53f8a054",
    79 => x"83bf5273",
    80 => x"70810555",
    81 => x"33517073",
    82 => x"70810555",
    83 => x"34ff1252",
    84 => x"718025eb",
    85 => x"38fbc053",
    86 => x"9f52a073",
    87 => x"70810555",
    88 => x"34ff1252",
    89 => x"718025f2",
    90 => x"38029005",
    91 => x"0d0402f4",
    92 => x"050d7453",
    93 => x"8e0bb0d4",
    94 => x"08258f38",
    95 => x"82b22db0",
    96 => x"d408ff05",
    97 => x"b0d40c82",
    98 => x"f404b0d4",
    99 => x"08b0d808",
   100 => x"5351728a",
   101 => x"2e098106",
   102 => x"b7387151",
   103 => x"719f24a0",
   104 => x"38b0d408",
   105 => x"a02911f8",
   106 => x"80115151",
   107 => x"a07134b0",
   108 => x"d8088105",
   109 => x"b0d80cb0",
   110 => x"d808519f",
   111 => x"7125e238",
   112 => x"800bb0d8",
   113 => x"0cb0d408",
   114 => x"8105b0d4",
   115 => x"0c83e404",
   116 => x"70a02912",
   117 => x"f8801151",
   118 => x"51727134",
   119 => x"b0d80881",
   120 => x"05b0d80c",
   121 => x"b0d808a0",
   122 => x"2e098106",
   123 => x"8e38800b",
   124 => x"b0d80cb0",
   125 => x"d4088105",
   126 => x"b0d40c02",
   127 => x"8c050d04",
   128 => x"02e8050d",
   129 => x"77795656",
   130 => x"880bfc16",
   131 => x"77712c8f",
   132 => x"06545254",
   133 => x"80537272",
   134 => x"25953871",
   135 => x"53fbe014",
   136 => x"51877134",
   137 => x"8114ff14",
   138 => x"545472f1",
   139 => x"387153f9",
   140 => x"1576712c",
   141 => x"87065351",
   142 => x"71802e8b",
   143 => x"38fbe014",
   144 => x"51717134",
   145 => x"81145472",
   146 => x"8e249538",
   147 => x"8f733153",
   148 => x"fbe01451",
   149 => x"a0713481",
   150 => x"14ff1454",
   151 => x"5472f138",
   152 => x"0298050d",
   153 => x"0402ec05",
   154 => x"0d800bb0",
   155 => x"e00cf68c",
   156 => x"08f69008",
   157 => x"71882c57",
   158 => x"5481ff06",
   159 => x"52747225",
   160 => x"88387155",
   161 => x"820bb0e0",
   162 => x"0c72882c",
   163 => x"7381ff06",
   164 => x"54547373",
   165 => x"258b3872",
   166 => x"b0e00884",
   167 => x"07b0e00c",
   168 => x"54b0dc08",
   169 => x"82055182",
   170 => x"0bb0dc0c",
   171 => x"830bf688",
   172 => x"0c74712b",
   173 => x"fecc0570",
   174 => x"9f2a1170",
   175 => x"812c7688",
   176 => x"29ff9405",
   177 => x"70812cb0",
   178 => x"e0085257",
   179 => x"52545151",
   180 => x"76802e85",
   181 => x"38708107",
   182 => x"5170f694",
   183 => x"0c710981",
   184 => x"05f6800c",
   185 => x"72098105",
   186 => x"f6840c02",
   187 => x"94050d04",
   188 => x"02f4050d",
   189 => x"74537270",
   190 => x"81055480",
   191 => x"f52d5271",
   192 => x"802e8938",
   193 => x"715182ee",
   194 => x"2d85f604",
   195 => x"028c050d",
   196 => x"040402f4",
   197 => x"050d7470",
   198 => x"8432b694",
   199 => x"0c708306",
   200 => x"525370ae",
   201 => x"d80b8805",
   202 => x"81b72d72",
   203 => x"892a7081",
   204 => x"06515170",
   205 => x"afa80b81",
   206 => x"b72d7283",
   207 => x"2a810673",
   208 => x"882a7081",
   209 => x"06515252",
   210 => x"70802e85",
   211 => x"38718207",
   212 => x"5271aef8",
   213 => x"0b81b72d",
   214 => x"72842c70",
   215 => x"83065151",
   216 => x"70af840b",
   217 => x"81b72d70",
   218 => x"b0c40c02",
   219 => x"8c050d04",
   220 => x"02f4050d",
   221 => x"b6940881",
   222 => x"c406afa8",
   223 => x"0b80f52d",
   224 => x"52527080",
   225 => x"2e863871",
   226 => x"84800752",
   227 => x"aee00b80",
   228 => x"f52d7207",
   229 => x"aef80b80",
   230 => x"f52d7081",
   231 => x"2a708106",
   232 => x"51535452",
   233 => x"70802e86",
   234 => x"38718280",
   235 => x"07527281",
   236 => x"06517080",
   237 => x"2e853871",
   238 => x"880752af",
   239 => x"840b80f5",
   240 => x"2d70842b",
   241 => x"73078432",
   242 => x"b0c40c51",
   243 => x"028c050d",
   244 => x"0402f805",
   245 => x"0da1842d",
   246 => x"80da51a2",
   247 => x"bb2db0c4",
   248 => x"08812a70",
   249 => x"81065152",
   250 => x"71802ee9",
   251 => x"38028805",
   252 => x"0d0402d4",
   253 => x"050d810b",
   254 => x"fec40c84",
   255 => x"b90bfec0",
   256 => x"0c840bfe",
   257 => x"c40ca0ec",
   258 => x"2da2ff2d",
   259 => x"a0d12da0",
   260 => x"d12d81f7",
   261 => x"2d815184",
   262 => x"e52da0d1",
   263 => x"2da0d12d",
   264 => x"815184e5",
   265 => x"2da9f851",
   266 => x"85f02d99",
   267 => x"8c2db0c4",
   268 => x"08802e82",
   269 => x"bc388bbf",
   270 => x"2db0c408",
   271 => x"53b0c408",
   272 => x"802e82b4",
   273 => x"389bc82d",
   274 => x"b0c40880",
   275 => x"2e8738aa",
   276 => x"905188e2",
   277 => x"0494d72d",
   278 => x"b0c40880",
   279 => x"2e8a38aa",
   280 => x"d05185f0",
   281 => x"2d87d12d",
   282 => x"ab985185",
   283 => x"f02dabb0",
   284 => x"52b0e451",
   285 => x"91db2db0",
   286 => x"c40881ff",
   287 => x"0653729d",
   288 => x"38abbc51",
   289 => x"85f02dab",
   290 => x"d452b0e4",
   291 => x"5191db2d",
   292 => x"b0c40881",
   293 => x"ff065372",
   294 => x"802e81cf",
   295 => x"38abe051",
   296 => x"85f02db0",
   297 => x"e8085780",
   298 => x"77595a76",
   299 => x"7a2e8b38",
   300 => x"811a7881",
   301 => x"2a595a77",
   302 => x"f738f71a",
   303 => x"5a807725",
   304 => x"80fe3879",
   305 => x"52775184",
   306 => x"802db0f0",
   307 => x"52b0e451",
   308 => x"94a02db0",
   309 => x"c40881ff",
   310 => x"06b0f05c",
   311 => x"53805972",
   312 => x"792e0981",
   313 => x"06b1388a",
   314 => x"aa047a70",
   315 => x"84055c08",
   316 => x"7081ff06",
   317 => x"71882c70",
   318 => x"81ff0673",
   319 => x"902c7081",
   320 => x"ff067598",
   321 => x"2afec80c",
   322 => x"fec80c58",
   323 => x"fec80c57",
   324 => x"fec80c84",
   325 => x"1a5a5376",
   326 => x"53848077",
   327 => x"25843884",
   328 => x"80537279",
   329 => x"24c4388a",
   330 => x"b004abfc",
   331 => x"5185f02d",
   332 => x"b0e45193",
   333 => x"f32dfc80",
   334 => x"17811959",
   335 => x"5789bd04",
   336 => x"820bfec4",
   337 => x"0c805184",
   338 => x"e52d0b0b",
   339 => x"0baea851",
   340 => x"a4a42d84",
   341 => x"b9518692",
   342 => x"2da1842d",
   343 => x"a4b42d86",
   344 => x"f02db0c4",
   345 => x"08fec00c",
   346 => x"8ad904ac",
   347 => x"905185f0",
   348 => x"2d820bfe",
   349 => x"c40c8053",
   350 => x"72b0c40c",
   351 => x"02ac050d",
   352 => x"0402e805",
   353 => x"0d77797b",
   354 => x"58555580",
   355 => x"53727625",
   356 => x"a3387470",
   357 => x"81055680",
   358 => x"f52d7470",
   359 => x"81055680",
   360 => x"f52d5252",
   361 => x"71712e86",
   362 => x"3881518b",
   363 => x"b6048113",
   364 => x"538b8d04",
   365 => x"805170b0",
   366 => x"c40c0298",
   367 => x"050d0402",
   368 => x"d8050d80",
   369 => x"0bb4f80c",
   370 => x"b0f05280",
   371 => x"519aa52d",
   372 => x"b0c40854",
   373 => x"b0c4088c",
   374 => x"38aca851",
   375 => x"85f02d73",
   376 => x"5590e404",
   377 => x"8056810b",
   378 => x"b59c0c88",
   379 => x"53acbc52",
   380 => x"b1a6518b",
   381 => x"812db0c4",
   382 => x"08762e09",
   383 => x"81068738",
   384 => x"b0c408b5",
   385 => x"9c0c8853",
   386 => x"acc852b1",
   387 => x"c2518b81",
   388 => x"2db0c408",
   389 => x"8738b0c4",
   390 => x"08b59c0c",
   391 => x"b59c0852",
   392 => x"acd4519d",
   393 => x"c22db59c",
   394 => x"08802e80",
   395 => x"f638b4b6",
   396 => x"0b80f52d",
   397 => x"b4b70b80",
   398 => x"f52d7198",
   399 => x"2b71902b",
   400 => x"07b4b80b",
   401 => x"80f52d70",
   402 => x"882b7207",
   403 => x"b4b90b80",
   404 => x"f52d7107",
   405 => x"b4ee0b80",
   406 => x"f52db4ef",
   407 => x"0b80f52d",
   408 => x"71882b07",
   409 => x"535f5452",
   410 => x"5a565755",
   411 => x"7381abaa",
   412 => x"2e098106",
   413 => x"8d387551",
   414 => x"9c972db0",
   415 => x"c408568d",
   416 => x"8f047382",
   417 => x"d4d52e87",
   418 => x"38acec51",
   419 => x"8dd004b0",
   420 => x"f0527551",
   421 => x"9aa52db0",
   422 => x"c40855b0",
   423 => x"c408802e",
   424 => x"83c23888",
   425 => x"53acc852",
   426 => x"b1c2518b",
   427 => x"812db0c4",
   428 => x"08893881",
   429 => x"0bb4f80c",
   430 => x"8dd60488",
   431 => x"53acbc52",
   432 => x"b1a6518b",
   433 => x"812db0c4",
   434 => x"08802e8a",
   435 => x"38ad8c51",
   436 => x"85f02d8e",
   437 => x"b004b4ee",
   438 => x"0b80f52d",
   439 => x"547380d5",
   440 => x"2e098106",
   441 => x"80ca38b4",
   442 => x"ef0b80f5",
   443 => x"2d547381",
   444 => x"aa2e0981",
   445 => x"06ba3880",
   446 => x"0bb0f00b",
   447 => x"80f52d56",
   448 => x"547481e9",
   449 => x"2e833881",
   450 => x"547481eb",
   451 => x"2e8c3880",
   452 => x"5573752e",
   453 => x"09810682",
   454 => x"cb38b0fb",
   455 => x"0b80f52d",
   456 => x"55748d38",
   457 => x"b0fc0b80",
   458 => x"f52d5473",
   459 => x"822e8638",
   460 => x"805590e4",
   461 => x"04b0fd0b",
   462 => x"80f52d70",
   463 => x"b4f00cff",
   464 => x"05b4f40c",
   465 => x"b0fe0b80",
   466 => x"f52db0ff",
   467 => x"0b80f52d",
   468 => x"58760577",
   469 => x"82802905",
   470 => x"70b4fc0c",
   471 => x"b1800b80",
   472 => x"f52d70b5",
   473 => x"900cb4f8",
   474 => x"08595758",
   475 => x"76802e81",
   476 => x"a3388853",
   477 => x"acc852b1",
   478 => x"c2518b81",
   479 => x"2db0c408",
   480 => x"81e238b4",
   481 => x"f0087084",
   482 => x"2bb5940c",
   483 => x"70b58c0c",
   484 => x"b1950b80",
   485 => x"f52db194",
   486 => x"0b80f52d",
   487 => x"71828029",
   488 => x"05b1960b",
   489 => x"80f52d70",
   490 => x"84808029",
   491 => x"12b1970b",
   492 => x"80f52d70",
   493 => x"81800a29",
   494 => x"1270b598",
   495 => x"0cb59008",
   496 => x"7129b4fc",
   497 => x"080570b5",
   498 => x"800cb19d",
   499 => x"0b80f52d",
   500 => x"b19c0b80",
   501 => x"f52d7182",
   502 => x"802905b1",
   503 => x"9e0b80f5",
   504 => x"2d708480",
   505 => x"802912b1",
   506 => x"9f0b80f5",
   507 => x"2d70982b",
   508 => x"81f00a06",
   509 => x"720570b5",
   510 => x"840cfe11",
   511 => x"7e297705",
   512 => x"b5880c52",
   513 => x"59524354",
   514 => x"5e515259",
   515 => x"525d5759",
   516 => x"5790e204",
   517 => x"b1820b80",
   518 => x"f52db181",
   519 => x"0b80f52d",
   520 => x"71828029",
   521 => x"0570b594",
   522 => x"0c70a029",
   523 => x"83ff0570",
   524 => x"892a70b5",
   525 => x"8c0cb187",
   526 => x"0b80f52d",
   527 => x"b1860b80",
   528 => x"f52d7182",
   529 => x"80290570",
   530 => x"b5980c7b",
   531 => x"71291e70",
   532 => x"b5880c7d",
   533 => x"b5840c73",
   534 => x"05b5800c",
   535 => x"555e5151",
   536 => x"55558155",
   537 => x"74b0c40c",
   538 => x"02a8050d",
   539 => x"0402ec05",
   540 => x"0d767087",
   541 => x"2c7180ff",
   542 => x"06555654",
   543 => x"b4f8088a",
   544 => x"3873882c",
   545 => x"7481ff06",
   546 => x"5455b0f0",
   547 => x"52b4fc08",
   548 => x"15519aa5",
   549 => x"2db0c408",
   550 => x"54b0c408",
   551 => x"802eb338",
   552 => x"b4f80880",
   553 => x"2e983872",
   554 => x"8429b0f0",
   555 => x"05700852",
   556 => x"539c972d",
   557 => x"b0c408f0",
   558 => x"0a065391",
   559 => x"d0047210",
   560 => x"b0f00570",
   561 => x"80e02d52",
   562 => x"539cc72d",
   563 => x"b0c40853",
   564 => x"725473b0",
   565 => x"c40c0294",
   566 => x"050d0402",
   567 => x"c8050d7f",
   568 => x"615f5b80",
   569 => x"0bb58408",
   570 => x"b5880859",
   571 => x"5d56b4f8",
   572 => x"08762e8a",
   573 => x"38b4f008",
   574 => x"842b5892",
   575 => x"8404b58c",
   576 => x"08842b58",
   577 => x"80597878",
   578 => x"2781a938",
   579 => x"788f06a0",
   580 => x"17575473",
   581 => x"8f38b0f0",
   582 => x"52765181",
   583 => x"17579aa5",
   584 => x"2db0f056",
   585 => x"807680f5",
   586 => x"2d565474",
   587 => x"742e8338",
   588 => x"81547481",
   589 => x"e52e80f6",
   590 => x"38817075",
   591 => x"06555d73",
   592 => x"802e80ea",
   593 => x"388b1680",
   594 => x"f52d9806",
   595 => x"5a7980de",
   596 => x"388b537d",
   597 => x"5275518b",
   598 => x"812db0c4",
   599 => x"0880cf38",
   600 => x"9c160851",
   601 => x"9c972db0",
   602 => x"c408841c",
   603 => x"0c9a1680",
   604 => x"e02d519c",
   605 => x"c72db0c4",
   606 => x"08b0c408",
   607 => x"881d0cb0",
   608 => x"c4085555",
   609 => x"b4f80880",
   610 => x"2e983894",
   611 => x"1680e02d",
   612 => x"519cc72d",
   613 => x"b0c40890",
   614 => x"2b83fff0",
   615 => x"0a067016",
   616 => x"51547388",
   617 => x"1c0c797b",
   618 => x"0c7c5493",
   619 => x"ea048119",
   620 => x"59928604",
   621 => x"b4f80880",
   622 => x"2eae387b",
   623 => x"5190ed2d",
   624 => x"b0c408b0",
   625 => x"c40880ff",
   626 => x"fffff806",
   627 => x"555c7380",
   628 => x"fffffff8",
   629 => x"2e9238b0",
   630 => x"c408fe05",
   631 => x"b4f00829",
   632 => x"b5800805",
   633 => x"57928404",
   634 => x"805473b0",
   635 => x"c40c02b8",
   636 => x"050d0402",
   637 => x"f4050d74",
   638 => x"70088105",
   639 => x"710c7008",
   640 => x"b4f40806",
   641 => x"5353718e",
   642 => x"38881308",
   643 => x"5190ed2d",
   644 => x"b0c40888",
   645 => x"140c810b",
   646 => x"b0c40c02",
   647 => x"8c050d04",
   648 => x"02f0050d",
   649 => x"75881108",
   650 => x"fe05b4f0",
   651 => x"0829b580",
   652 => x"08117208",
   653 => x"b4f40806",
   654 => x"05795553",
   655 => x"54549aa5",
   656 => x"2db0c408",
   657 => x"53b0c408",
   658 => x"802e8338",
   659 => x"815372b0",
   660 => x"c40c0290",
   661 => x"050d04b4",
   662 => x"f808b0c4",
   663 => x"0c0402f4",
   664 => x"050dd452",
   665 => x"81ff720c",
   666 => x"71085381",
   667 => x"ff720c72",
   668 => x"882b83fe",
   669 => x"80067208",
   670 => x"7081ff06",
   671 => x"51525381",
   672 => x"ff720c72",
   673 => x"7107882b",
   674 => x"72087081",
   675 => x"ff065152",
   676 => x"5381ff72",
   677 => x"0c727107",
   678 => x"882b7208",
   679 => x"7081ff06",
   680 => x"7207b0c4",
   681 => x"0c525302",
   682 => x"8c050d04",
   683 => x"02f4050d",
   684 => x"74767181",
   685 => x"ff06d40c",
   686 => x"5353b5a0",
   687 => x"08853871",
   688 => x"892b5271",
   689 => x"982ad40c",
   690 => x"71902a70",
   691 => x"81ff06d4",
   692 => x"0c517188",
   693 => x"2a7081ff",
   694 => x"06d40c51",
   695 => x"7181ff06",
   696 => x"d40c7290",
   697 => x"2a7081ff",
   698 => x"06d40c51",
   699 => x"d4087081",
   700 => x"ff065151",
   701 => x"82b8bf52",
   702 => x"7081ff2e",
   703 => x"09810694",
   704 => x"3881ff0b",
   705 => x"d40cd408",
   706 => x"7081ff06",
   707 => x"ff145451",
   708 => x"5171e538",
   709 => x"70b0c40c",
   710 => x"028c050d",
   711 => x"0402fc05",
   712 => x"0d81c751",
   713 => x"81ff0bd4",
   714 => x"0cff1151",
   715 => x"708025f4",
   716 => x"38028405",
   717 => x"0d0402f0",
   718 => x"050d969d",
   719 => x"2d819c9f",
   720 => x"53805287",
   721 => x"fc80f751",
   722 => x"95ac2db0",
   723 => x"c40854b0",
   724 => x"c408812e",
   725 => x"098106a3",
   726 => x"3881ff0b",
   727 => x"d40c820a",
   728 => x"52849c80",
   729 => x"e95195ac",
   730 => x"2db0c408",
   731 => x"8b3881ff",
   732 => x"0bd40c73",
   733 => x"53978104",
   734 => x"969d2dff",
   735 => x"135372c1",
   736 => x"3872b0c4",
   737 => x"0c029005",
   738 => x"0d0402f4",
   739 => x"050d81ff",
   740 => x"0bd40c93",
   741 => x"53805287",
   742 => x"fc80c151",
   743 => x"95ac2db0",
   744 => x"c4088b38",
   745 => x"81ff0bd4",
   746 => x"0c815397",
   747 => x"b704969d",
   748 => x"2dff1353",
   749 => x"72df3872",
   750 => x"b0c40c02",
   751 => x"8c050d04",
   752 => x"02f0050d",
   753 => x"969d2d83",
   754 => x"aa52849c",
   755 => x"80c85195",
   756 => x"ac2db0c4",
   757 => x"08812e09",
   758 => x"81069238",
   759 => x"94de2db0",
   760 => x"c40883ff",
   761 => x"ff065372",
   762 => x"83aa2e97",
   763 => x"38978a2d",
   764 => x"97fe0481",
   765 => x"54998304",
   766 => x"adac5185",
   767 => x"f02d8054",
   768 => x"99830481",
   769 => x"ff0bd40c",
   770 => x"b15396b6",
   771 => x"2db0c408",
   772 => x"802e80e0",
   773 => x"38805287",
   774 => x"fc80fa51",
   775 => x"95ac2db0",
   776 => x"c40880c6",
   777 => x"38b0c408",
   778 => x"52adc851",
   779 => x"9dc22d81",
   780 => x"ff0bd40c",
   781 => x"d4087081",
   782 => x"ff067054",
   783 => x"add45351",
   784 => x"539dc22d",
   785 => x"81ff0bd4",
   786 => x"0c81ff0b",
   787 => x"d40c81ff",
   788 => x"0bd40c81",
   789 => x"ff0bd40c",
   790 => x"72862a70",
   791 => x"81067056",
   792 => x"51537280",
   793 => x"2e9d3897",
   794 => x"f304b0c4",
   795 => x"0852adc8",
   796 => x"519dc22d",
   797 => x"72822efe",
   798 => x"ff38ff13",
   799 => x"5372ff8a",
   800 => x"38725473",
   801 => x"b0c40c02",
   802 => x"90050d04",
   803 => x"02f4050d",
   804 => x"810bb5a0",
   805 => x"0cd00870",
   806 => x"8f2a7081",
   807 => x"06515153",
   808 => x"72f33872",
   809 => x"d00c969d",
   810 => x"2dd00870",
   811 => x"8f2a7081",
   812 => x"06515153",
   813 => x"72f33881",
   814 => x"0bd00c87",
   815 => x"53805284",
   816 => x"d480c051",
   817 => x"95ac2db0",
   818 => x"c408812e",
   819 => x"9a387282",
   820 => x"2e098106",
   821 => x"8c38ade4",
   822 => x"5185f02d",
   823 => x"80539a9c",
   824 => x"04ff1353",
   825 => x"72d73897",
   826 => x"c02db0c4",
   827 => x"08b5a00c",
   828 => x"b0c4088b",
   829 => x"38815287",
   830 => x"fc80d051",
   831 => x"95ac2d81",
   832 => x"ff0bd40c",
   833 => x"d008708f",
   834 => x"2a708106",
   835 => x"51515372",
   836 => x"f33872d0",
   837 => x"0c81ff0b",
   838 => x"d40c8153",
   839 => x"72b0c40c",
   840 => x"028c050d",
   841 => x"0402e005",
   842 => x"0d797b57",
   843 => x"57805881",
   844 => x"ff0bd40c",
   845 => x"d008708f",
   846 => x"2a708106",
   847 => x"51515473",
   848 => x"f3388281",
   849 => x"0bd00c81",
   850 => x"ff0bd40c",
   851 => x"765287fc",
   852 => x"80d15195",
   853 => x"ac2d80db",
   854 => x"c6df55b0",
   855 => x"c408802e",
   856 => x"9038b0c4",
   857 => x"08537652",
   858 => x"adfc519d",
   859 => x"c22d9bbf",
   860 => x"0481ff0b",
   861 => x"d40cd408",
   862 => x"7081ff06",
   863 => x"51547381",
   864 => x"fe2e0981",
   865 => x"069d3880",
   866 => x"ff5494de",
   867 => x"2db0c408",
   868 => x"76708405",
   869 => x"580cff14",
   870 => x"54738025",
   871 => x"ed388158",
   872 => x"9ba904ff",
   873 => x"155574c9",
   874 => x"3881ff0b",
   875 => x"d40cd008",
   876 => x"708f2a70",
   877 => x"81065151",
   878 => x"5473f338",
   879 => x"73d00c77",
   880 => x"b0c40c02",
   881 => x"a0050d04",
   882 => x"b5a008b0",
   883 => x"c40c0402",
   884 => x"e8050d80",
   885 => x"78575575",
   886 => x"70840557",
   887 => x"08538054",
   888 => x"72982a73",
   889 => x"882b5452",
   890 => x"71802ea2",
   891 => x"38c00870",
   892 => x"882a7081",
   893 => x"06515151",
   894 => x"70802ef1",
   895 => x"3871c00c",
   896 => x"81158115",
   897 => x"55558374",
   898 => x"25d63871",
   899 => x"ca3874b0",
   900 => x"c40c0298",
   901 => x"050d0402",
   902 => x"f4050d74",
   903 => x"70882a83",
   904 => x"fe800670",
   905 => x"72982a07",
   906 => x"72882b87",
   907 => x"fc808006",
   908 => x"73982b81",
   909 => x"f00a0671",
   910 => x"730707b0",
   911 => x"c40c5651",
   912 => x"5351028c",
   913 => x"050d0402",
   914 => x"f8050d02",
   915 => x"8e0580f5",
   916 => x"2d74882b",
   917 => x"077083ff",
   918 => x"ff06b0c4",
   919 => x"0c510288",
   920 => x"050d0402",
   921 => x"ec050d76",
   922 => x"53805572",
   923 => x"75258b38",
   924 => x"ad5182ee",
   925 => x"2d720981",
   926 => x"05537280",
   927 => x"2eb53887",
   928 => x"54729c2a",
   929 => x"73842b54",
   930 => x"5271802e",
   931 => x"83388155",
   932 => x"89722587",
   933 => x"38b71252",
   934 => x"9d9e04b0",
   935 => x"12527480",
   936 => x"2e863871",
   937 => x"5182ee2d",
   938 => x"ff145473",
   939 => x"8025d238",
   940 => x"9db804b0",
   941 => x"5182ee2d",
   942 => x"800bb0c4",
   943 => x"0c029405",
   944 => x"0d0402c0",
   945 => x"050d0280",
   946 => x"c4055780",
   947 => x"70787084",
   948 => x"055a0872",
   949 => x"415f5d58",
   950 => x"7c708405",
   951 => x"5e085a80",
   952 => x"5b79982a",
   953 => x"7a882b5b",
   954 => x"56758638",
   955 => x"775f9fba",
   956 => x"047d802e",
   957 => x"81a23880",
   958 => x"5e7580e4",
   959 => x"2e8a3875",
   960 => x"80f82e09",
   961 => x"81068938",
   962 => x"76841871",
   963 => x"085e5854",
   964 => x"7580e42e",
   965 => x"9f387580",
   966 => x"e4268a38",
   967 => x"7580e32e",
   968 => x"be389eea",
   969 => x"047580f3",
   970 => x"2ea33875",
   971 => x"80f82e89",
   972 => x"389eea04",
   973 => x"8a539ebb",
   974 => x"049053b5",
   975 => x"a4527b51",
   976 => x"9ce32db0",
   977 => x"c408b5a4",
   978 => x"5a559efa",
   979 => x"04768418",
   980 => x"71087054",
   981 => x"5b58549b",
   982 => x"cf2d8055",
   983 => x"9efa0476",
   984 => x"84187108",
   985 => x"5858549f",
   986 => x"a504a551",
   987 => x"82ee2d75",
   988 => x"5182ee2d",
   989 => x"8218589f",
   990 => x"ad0474ff",
   991 => x"16565480",
   992 => x"7425aa38",
   993 => x"78708105",
   994 => x"5a80f52d",
   995 => x"70525682",
   996 => x"ee2d8118",
   997 => x"589efa04",
   998 => x"75a52e09",
   999 => x"81068638",
  1000 => x"815e9fad",
  1001 => x"04755182",
  1002 => x"ee2d8118",
  1003 => x"58811b5b",
  1004 => x"837b25fe",
  1005 => x"ac3875fe",
  1006 => x"9f387eb0",
  1007 => x"c40c0280",
  1008 => x"c0050d04",
  1009 => x"02fc050d",
  1010 => x"72518071",
  1011 => x"0c800b84",
  1012 => x"120c0284",
  1013 => x"050d0402",
  1014 => x"f0050d75",
  1015 => x"70088412",
  1016 => x"08535353",
  1017 => x"ff547171",
  1018 => x"2e9b3884",
  1019 => x"13087084",
  1020 => x"29148b11",
  1021 => x"80f52d84",
  1022 => x"16088111",
  1023 => x"87068418",
  1024 => x"0c525651",
  1025 => x"5173b0c4",
  1026 => x"0c029005",
  1027 => x"0d0402f8",
  1028 => x"050da385",
  1029 => x"2de00870",
  1030 => x"8b2a7081",
  1031 => x"06515252",
  1032 => x"70802e9d",
  1033 => x"38b5e408",
  1034 => x"708429b5",
  1035 => x"ec057381",
  1036 => x"ff06710c",
  1037 => x"5151b5e4",
  1038 => x"08811187",
  1039 => x"06b5e40c",
  1040 => x"51800bb6",
  1041 => x"8c0ca2f8",
  1042 => x"2da2ff2d",
  1043 => x"0288050d",
  1044 => x"0402fc05",
  1045 => x"0da3852d",
  1046 => x"810bb68c",
  1047 => x"0ca2ff2d",
  1048 => x"b68c0851",
  1049 => x"70fa3802",
  1050 => x"84050d04",
  1051 => x"02fc050d",
  1052 => x"b5e4519f",
  1053 => x"c42da08e",
  1054 => x"51a2f42d",
  1055 => x"a29e2d02",
  1056 => x"84050d04",
  1057 => x"02f4050d",
  1058 => x"a28604b0",
  1059 => x"c40881f0",
  1060 => x"2e098106",
  1061 => x"8938810b",
  1062 => x"b0b80ca2",
  1063 => x"8604b0c4",
  1064 => x"0881e02e",
  1065 => x"09810689",
  1066 => x"38810bb0",
  1067 => x"bc0ca286",
  1068 => x"04b0c408",
  1069 => x"52b0bc08",
  1070 => x"802e8838",
  1071 => x"b0c40881",
  1072 => x"80055271",
  1073 => x"842c728f",
  1074 => x"065353b0",
  1075 => x"b808802e",
  1076 => x"99387284",
  1077 => x"29aff805",
  1078 => x"72138171",
  1079 => x"2b700973",
  1080 => x"0806730c",
  1081 => x"515353a1",
  1082 => x"fc047284",
  1083 => x"29aff805",
  1084 => x"72138371",
  1085 => x"2b720807",
  1086 => x"720c5353",
  1087 => x"800bb0bc",
  1088 => x"0c800bb0",
  1089 => x"b80cb5e4",
  1090 => x"519fd72d",
  1091 => x"b0c408ff",
  1092 => x"24fef838",
  1093 => x"800bb0c4",
  1094 => x"0c028c05",
  1095 => x"0d0402f8",
  1096 => x"050daff8",
  1097 => x"528f5180",
  1098 => x"72708405",
  1099 => x"540cff11",
  1100 => x"51708025",
  1101 => x"f2380288",
  1102 => x"050d0402",
  1103 => x"f0050d75",
  1104 => x"51a3852d",
  1105 => x"70822cfc",
  1106 => x"06aff811",
  1107 => x"72109e06",
  1108 => x"71087072",
  1109 => x"2a708306",
  1110 => x"82742b70",
  1111 => x"09740676",
  1112 => x"0c545156",
  1113 => x"57535153",
  1114 => x"a2ff2d71",
  1115 => x"b0c40c02",
  1116 => x"90050d04",
  1117 => x"71980c04",
  1118 => x"ffb008b0",
  1119 => x"c40c0481",
  1120 => x"0bffb00c",
  1121 => x"04800bff",
  1122 => x"b00c0402",
  1123 => x"fc050d80",
  1124 => x"0bb0c00c",
  1125 => x"805184e5",
  1126 => x"2d028405",
  1127 => x"0d0402f0",
  1128 => x"050db690",
  1129 => x"085481f7",
  1130 => x"2d800bb6",
  1131 => x"980c7308",
  1132 => x"802e80eb",
  1133 => x"38820bb0",
  1134 => x"d80cb698",
  1135 => x"088f06b0",
  1136 => x"d40c7308",
  1137 => x"5271812e",
  1138 => x"a4387183",
  1139 => x"2e098106",
  1140 => x"b9388814",
  1141 => x"80f52d84",
  1142 => x"1508ae9c",
  1143 => x"53545285",
  1144 => x"f02d7184",
  1145 => x"29137008",
  1146 => x"5252a48e",
  1147 => x"04b69408",
  1148 => x"8815082c",
  1149 => x"70810651",
  1150 => x"5271802e",
  1151 => x"8738aea0",
  1152 => x"51a48704",
  1153 => x"aea45185",
  1154 => x"f02d8414",
  1155 => x"085185f0",
  1156 => x"2db69808",
  1157 => x"8105b698",
  1158 => x"0c8c1454",
  1159 => x"a3ae0402",
  1160 => x"90050d04",
  1161 => x"71b6900c",
  1162 => x"a39e2db6",
  1163 => x"9808ff05",
  1164 => x"b69c0c04",
  1165 => x"02f0050d",
  1166 => x"8751a2bb",
  1167 => x"2db0c408",
  1168 => x"812a7081",
  1169 => x"06515271",
  1170 => x"802e8e38",
  1171 => x"b0c00881",
  1172 => x"3270b0c0",
  1173 => x"0c5184e5",
  1174 => x"2db0c008",
  1175 => x"963880da",
  1176 => x"51a2bb2d",
  1177 => x"81f551a2",
  1178 => x"bb2d81f2",
  1179 => x"51a2bb2d",
  1180 => x"a78c0481",
  1181 => x"f551a2bb",
  1182 => x"2db0c408",
  1183 => x"812a7081",
  1184 => x"06515271",
  1185 => x"802e8f38",
  1186 => x"b69c0852",
  1187 => x"71802e86",
  1188 => x"38ff12b6",
  1189 => x"9c0c81f2",
  1190 => x"51a2bb2d",
  1191 => x"b0c40881",
  1192 => x"2a708106",
  1193 => x"51527180",
  1194 => x"2e9538b6",
  1195 => x"9808ff05",
  1196 => x"b69c0854",
  1197 => x"52727225",
  1198 => x"86388113",
  1199 => x"b69c0c80",
  1200 => x"da51a2bb",
  1201 => x"2db0c408",
  1202 => x"812a7081",
  1203 => x"06515271",
  1204 => x"802e80fb",
  1205 => x"38b69008",
  1206 => x"b69c0855",
  1207 => x"5373802e",
  1208 => x"8a388c13",
  1209 => x"ff155553",
  1210 => x"a5dd0472",
  1211 => x"08527182",
  1212 => x"2ea63871",
  1213 => x"82268938",
  1214 => x"71812ea5",
  1215 => x"38a6cf04",
  1216 => x"71832ead",
  1217 => x"3871842e",
  1218 => x"09810680",
  1219 => x"c2388813",
  1220 => x"0851a4a4",
  1221 => x"2da6cf04",
  1222 => x"88130852",
  1223 => x"712da6cf",
  1224 => x"04810b88",
  1225 => x"14082bb6",
  1226 => x"940832b6",
  1227 => x"940ca6cc",
  1228 => x"04881380",
  1229 => x"f52d8105",
  1230 => x"8b1480f5",
  1231 => x"2d535471",
  1232 => x"74248338",
  1233 => x"80547388",
  1234 => x"1481b72d",
  1235 => x"a39e2d80",
  1236 => x"54800bb0",
  1237 => x"d80c738f",
  1238 => x"06b0d40c",
  1239 => x"a05273b6",
  1240 => x"9c082e09",
  1241 => x"81069838",
  1242 => x"b69808ff",
  1243 => x"05743270",
  1244 => x"09810570",
  1245 => x"72079f2a",
  1246 => x"91713151",
  1247 => x"51535371",
  1248 => x"5182ee2d",
  1249 => x"8114548e",
  1250 => x"7425c638",
  1251 => x"0290050d",
  1252 => x"04000000",
  1253 => x"00ffffff",
  1254 => x"ff00ffff",
  1255 => x"ffff00ff",
  1256 => x"ffffff00",
  1257 => x"44495020",
  1258 => x"53776974",
  1259 => x"63686573",
  1260 => x"20100000",
  1261 => x"52657365",
  1262 => x"74000000",
  1263 => x"45786974",
  1264 => x"00000000",
  1265 => x"53442043",
  1266 => x"61726400",
  1267 => x"4a617061",
  1268 => x"6e657365",
  1269 => x"206b6579",
  1270 => x"626f6172",
  1271 => x"64206c61",
  1272 => x"796f7574",
  1273 => x"00000000",
  1274 => x"54757262",
  1275 => x"6f202831",
  1276 => x"302e3734",
  1277 => x"4d487a29",
  1278 => x"00000000",
  1279 => x"4261636b",
  1280 => x"00000000",
  1281 => x"32303438",
  1282 => x"4c422052",
  1283 => x"414d0000",
  1284 => x"34303936",
  1285 => x"4b422052",
  1286 => x"414d0000",
  1287 => x"536c323a",
  1288 => x"204e6f6e",
  1289 => x"65000000",
  1290 => x"536c323a",
  1291 => x"20455345",
  1292 => x"2d534343",
  1293 => x"20314d42",
  1294 => x"2f534343",
  1295 => x"2d490000",
  1296 => x"536c323a",
  1297 => x"20455345",
  1298 => x"2d52414d",
  1299 => x"20314d42",
  1300 => x"2f415343",
  1301 => x"49493800",
  1302 => x"536c323a",
  1303 => x"20455345",
  1304 => x"2d52414d",
  1305 => x"20314d42",
  1306 => x"2f415343",
  1307 => x"49493136",
  1308 => x"00000000",
  1309 => x"536c313a",
  1310 => x"204e6f6e",
  1311 => x"65000000",
  1312 => x"536c313a",
  1313 => x"20455345",
  1314 => x"2d534343",
  1315 => x"20314d42",
  1316 => x"2f534343",
  1317 => x"2d490000",
  1318 => x"536c313a",
  1319 => x"204d6567",
  1320 => x"6152414d",
  1321 => x"00000000",
  1322 => x"56474120",
  1323 => x"2d203331",
  1324 => x"4b487a2c",
  1325 => x"20363048",
  1326 => x"7a000000",
  1327 => x"56474120",
  1328 => x"2d203331",
  1329 => x"4b487a2c",
  1330 => x"20353048",
  1331 => x"7a000000",
  1332 => x"53434152",
  1333 => x"54202d20",
  1334 => x"31354b48",
  1335 => x"7a2c2035",
  1336 => x"30487a20",
  1337 => x"52474200",
  1338 => x"54562f53",
  1339 => x"6f756e64",
  1340 => x"202d2031",
  1341 => x"35487a00",
  1342 => x"496e6974",
  1343 => x"69616c69",
  1344 => x"7a696e67",
  1345 => x"20534420",
  1346 => x"63617264",
  1347 => x"0a000000",
  1348 => x"53444843",
  1349 => x"20636172",
  1350 => x"64206465",
  1351 => x"74656374",
  1352 => x"65642062",
  1353 => x"7574206e",
  1354 => x"6f740a73",
  1355 => x"7570706f",
  1356 => x"72746564",
  1357 => x"202d2064",
  1358 => x"69736162",
  1359 => x"6c696e67",
  1360 => x"20534420",
  1361 => x"63617264",
  1362 => x"0a10204f",
  1363 => x"4b0a0000",
  1364 => x"46617433",
  1365 => x"32206669",
  1366 => x"6c657379",
  1367 => x"7374656d",
  1368 => x"20646574",
  1369 => x"65637465",
  1370 => x"64206275",
  1371 => x"74206e6f",
  1372 => x"740a7375",
  1373 => x"70706f72",
  1374 => x"74656420",
  1375 => x"2d206469",
  1376 => x"7361626c",
  1377 => x"696e6720",
  1378 => x"53442063",
  1379 => x"6172640a",
  1380 => x"10204f4b",
  1381 => x"0a000000",
  1382 => x"54727969",
  1383 => x"6e67204d",
  1384 => x"53583342",
  1385 => x"494f532e",
  1386 => x"5359532e",
  1387 => x"2e2e0a00",
  1388 => x"4d535833",
  1389 => x"42494f53",
  1390 => x"53595300",
  1391 => x"54727969",
  1392 => x"6e672042",
  1393 => x"494f535f",
  1394 => x"4d32502e",
  1395 => x"524f4d2e",
  1396 => x"2e2e0a00",
  1397 => x"42494f53",
  1398 => x"5f4d3250",
  1399 => x"524f4d00",
  1400 => x"4f70656e",
  1401 => x"65642042",
  1402 => x"494f532c",
  1403 => x"206c6f61",
  1404 => x"64696e67",
  1405 => x"2e2e2e0a",
  1406 => x"00000000",
  1407 => x"52656164",
  1408 => x"20626c6f",
  1409 => x"636b2066",
  1410 => x"61696c65",
  1411 => x"640a0000",
  1412 => x"4c6f6164",
  1413 => x"696e6720",
  1414 => x"42494f53",
  1415 => x"20666169",
  1416 => x"6c65640a",
  1417 => x"00000000",
  1418 => x"52656164",
  1419 => x"206f6620",
  1420 => x"4d425220",
  1421 => x"6661696c",
  1422 => x"65640a00",
  1423 => x"46415431",
  1424 => x"36202020",
  1425 => x"00000000",
  1426 => x"46415433",
  1427 => x"32202020",
  1428 => x"00000000",
  1429 => x"25642070",
  1430 => x"61727469",
  1431 => x"74696f6e",
  1432 => x"7320666f",
  1433 => x"756e640a",
  1434 => x"00000000",
  1435 => x"4e6f2070",
  1436 => x"61727469",
  1437 => x"74696f6e",
  1438 => x"20736967",
  1439 => x"6e617475",
  1440 => x"72652066",
  1441 => x"6f756e64",
  1442 => x"0a000000",
  1443 => x"556e7375",
  1444 => x"70706f72",
  1445 => x"74656420",
  1446 => x"70617274",
  1447 => x"6974696f",
  1448 => x"6e207479",
  1449 => x"7065210a",
  1450 => x"00000000",
  1451 => x"53444843",
  1452 => x"20496e69",
  1453 => x"7469616c",
  1454 => x"697a6174",
  1455 => x"696f6e20",
  1456 => x"6572726f",
  1457 => x"72210a00",
  1458 => x"434d4435",
  1459 => x"38202564",
  1460 => x"0a202000",
  1461 => x"434d4435",
  1462 => x"385f3220",
  1463 => x"25640a20",
  1464 => x"20000000",
  1465 => x"53442063",
  1466 => x"61726420",
  1467 => x"72657365",
  1468 => x"74206661",
  1469 => x"696c6564",
  1470 => x"210a0000",
  1471 => x"52656164",
  1472 => x"20636f6d",
  1473 => x"6d616e64",
  1474 => x"20666169",
  1475 => x"6c656420",
  1476 => x"61742025",
  1477 => x"64202825",
  1478 => x"64290a00",
  1479 => x"16200000",
  1480 => x"14200000",
  1481 => x"15200000",
  1482 => x"00000004",
  1483 => x"000013a4",
  1484 => x"00001758",
  1485 => x"00000002",
  1486 => x"000013b4",
  1487 => x"00000311",
  1488 => x"00000002",
  1489 => x"000013bc",
  1490 => x"0000118b",
  1491 => x"00000000",
  1492 => x"00000000",
  1493 => x"00000000",
  1494 => x"00000003",
  1495 => x"000017e8",
  1496 => x"00000004",
  1497 => x"00000001",
  1498 => x"000013c4",
  1499 => x"00000002",
  1500 => x"00000003",
  1501 => x"000017dc",
  1502 => x"00000003",
  1503 => x"00000003",
  1504 => x"000017cc",
  1505 => x"00000004",
  1506 => x"00000001",
  1507 => x"000013cc",
  1508 => x"00000006",
  1509 => x"00000001",
  1510 => x"000013e8",
  1511 => x"00000007",
  1512 => x"00000003",
  1513 => x"000017c4",
  1514 => x"00000002",
  1515 => x"00000004",
  1516 => x"000013fc",
  1517 => x"00001728",
  1518 => x"00000000",
  1519 => x"00000000",
  1520 => x"00000000",
  1521 => x"00001404",
  1522 => x"00001410",
  1523 => x"0000141c",
  1524 => x"00001428",
  1525 => x"00001440",
  1526 => x"00001458",
  1527 => x"00001474",
  1528 => x"00001480",
  1529 => x"00001498",
  1530 => x"000014a8",
  1531 => x"000014bc",
  1532 => x"000014d0",
  1533 => x"000014e8",
  1534 => x"00000000",
  1535 => x"00000000",
  1536 => x"00000000",
  1537 => x"00000000",
  1538 => x"00000000",
  1539 => x"00000000",
  1540 => x"00000000",
  1541 => x"00000000",
  1542 => x"00000000",
  1543 => x"00000000",
  1544 => x"00000000",
  1545 => x"00000000",
  1546 => x"00000000",
  1547 => x"00000000",
  1548 => x"00000000",
  1549 => x"00000000",
  1550 => x"00000000",
  1551 => x"00000000",
  1552 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

