-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"000b0b0b",
     4 => x"0b8c04ff",
     5 => x"0d800404",
     6 => x"00000017",
     7 => x"00000000",
     8 => x"0b0b0bb7",
     9 => x"f8080b0b",
    10 => x"0bb7fc08",
    11 => x"0b0b0bb8",
    12 => x"80080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"b8800c0b",
    16 => x"0b0bb7fc",
    17 => x"0c0b0b0b",
    18 => x"b7f80c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0baed8",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"b7f870bd",
    57 => x"b0278b38",
    58 => x"80717084",
    59 => x"05530c81",
    60 => x"e2048c51",
    61 => x"8d9b0402",
    62 => x"fc050df8",
    63 => x"80518f0b",
    64 => x"b8880c9f",
    65 => x"0bb88c0c",
    66 => x"a0717081",
    67 => x"055334b8",
    68 => x"8c08ff05",
    69 => x"b88c0cb8",
    70 => x"8c088025",
    71 => x"eb38b888",
    72 => x"08ff05b8",
    73 => x"880cb888",
    74 => x"088025d7",
    75 => x"38028405",
    76 => x"0d0402f0",
    77 => x"050df880",
    78 => x"53f8a054",
    79 => x"83bf5273",
    80 => x"70810555",
    81 => x"33517073",
    82 => x"70810555",
    83 => x"34ff1252",
    84 => x"718025eb",
    85 => x"38fbc053",
    86 => x"9f52a073",
    87 => x"70810555",
    88 => x"34ff1252",
    89 => x"718025f2",
    90 => x"38029005",
    91 => x"0d0402f4",
    92 => x"050d7453",
    93 => x"8e0bb888",
    94 => x"08258f38",
    95 => x"82b22db8",
    96 => x"8808ff05",
    97 => x"b8880c82",
    98 => x"f404b888",
    99 => x"08b88c08",
   100 => x"5351728a",
   101 => x"2e098106",
   102 => x"b7387151",
   103 => x"719f24a0",
   104 => x"38b88808",
   105 => x"a02911f8",
   106 => x"80115151",
   107 => x"a07134b8",
   108 => x"8c088105",
   109 => x"b88c0cb8",
   110 => x"8c08519f",
   111 => x"7125e238",
   112 => x"800bb88c",
   113 => x"0cb88808",
   114 => x"8105b888",
   115 => x"0c83e404",
   116 => x"70a02912",
   117 => x"f8801151",
   118 => x"51727134",
   119 => x"b88c0881",
   120 => x"05b88c0c",
   121 => x"b88c08a0",
   122 => x"2e098106",
   123 => x"8e38800b",
   124 => x"b88c0cb8",
   125 => x"88088105",
   126 => x"b8880c02",
   127 => x"8c050d04",
   128 => x"02e8050d",
   129 => x"77795656",
   130 => x"880bfc16",
   131 => x"77712c8f",
   132 => x"06545254",
   133 => x"80537272",
   134 => x"25953871",
   135 => x"53fbe014",
   136 => x"51877134",
   137 => x"8114ff14",
   138 => x"545472f1",
   139 => x"387153f9",
   140 => x"1576712c",
   141 => x"87065351",
   142 => x"71802e8b",
   143 => x"38fbe014",
   144 => x"51717134",
   145 => x"81145472",
   146 => x"8e249538",
   147 => x"8f733153",
   148 => x"fbe01451",
   149 => x"a0713481",
   150 => x"14ff1454",
   151 => x"5472f138",
   152 => x"0298050d",
   153 => x"0402ec05",
   154 => x"0d800bb8",
   155 => x"900cf68c",
   156 => x"08f69008",
   157 => x"71882c56",
   158 => x"5481ff06",
   159 => x"52737225",
   160 => x"88387154",
   161 => x"820bb890",
   162 => x"0c72882c",
   163 => x"7381ff06",
   164 => x"54557473",
   165 => x"258b3872",
   166 => x"b8900884",
   167 => x"07b8900c",
   168 => x"5573842b",
   169 => x"86a07125",
   170 => x"83713170",
   171 => x"0b0b0bb4",
   172 => x"d80c8171",
   173 => x"2bff05f6",
   174 => x"880cfecc",
   175 => x"13ff122c",
   176 => x"788829ff",
   177 => x"94057081",
   178 => x"2cb89008",
   179 => x"52585255",
   180 => x"51525476",
   181 => x"802e8538",
   182 => x"70810751",
   183 => x"70f6940c",
   184 => x"71098105",
   185 => x"f6800c72",
   186 => x"098105f6",
   187 => x"840c0294",
   188 => x"050d0402",
   189 => x"f4050d74",
   190 => x"53727081",
   191 => x"055480f5",
   192 => x"2d527180",
   193 => x"2e893871",
   194 => x"5182ee2d",
   195 => x"85f90402",
   196 => x"8c050d04",
   197 => x"02f8050d",
   198 => x"a6902d80",
   199 => x"da51a7c7",
   200 => x"2db7f808",
   201 => x"812a7081",
   202 => x"06515271",
   203 => x"802ee938",
   204 => x"0288050d",
   205 => x"0402f405",
   206 => x"0dbda008",
   207 => x"99c406b6",
   208 => x"d40b80f5",
   209 => x"2d525270",
   210 => x"802e8638",
   211 => x"71848007",
   212 => x"52b68c0b",
   213 => x"80f52d72",
   214 => x"07b6b00b",
   215 => x"80f52d70",
   216 => x"812a7081",
   217 => x"06515354",
   218 => x"5270802e",
   219 => x"86387182",
   220 => x"80075272",
   221 => x"81065170",
   222 => x"802e8538",
   223 => x"71880752",
   224 => x"b6bc0b80",
   225 => x"f52d7084",
   226 => x"2b730781",
   227 => x"8432b7f8",
   228 => x"0c51028c",
   229 => x"050d0402",
   230 => x"f4050d74",
   231 => x"70818432",
   232 => x"bda00c70",
   233 => x"83065253",
   234 => x"70b6840b",
   235 => x"880581b7",
   236 => x"2d72892a",
   237 => x"70810651",
   238 => x"5170b6d4",
   239 => x"0b81b72d",
   240 => x"72832a81",
   241 => x"0673882a",
   242 => x"70810651",
   243 => x"52527080",
   244 => x"2e853871",
   245 => x"82075271",
   246 => x"b6b00b81",
   247 => x"b72d7284",
   248 => x"2c708306",
   249 => x"515170b6",
   250 => x"bc0b81b7",
   251 => x"2d70b7f8",
   252 => x"0c028c05",
   253 => x"0d0402f4",
   254 => x"050db5bc",
   255 => x"0b881180",
   256 => x"f52d8c12",
   257 => x"881180f5",
   258 => x"2d70842b",
   259 => x"73078c13",
   260 => x"881180f5",
   261 => x"2d70882b",
   262 => x"73079413",
   263 => x"80f52d70",
   264 => x"8c2b7207",
   265 => x"b7f80c53",
   266 => x"53535353",
   267 => x"56525351",
   268 => x"028c050d",
   269 => x"0402f405",
   270 => x"0d74b5bc",
   271 => x"71870655",
   272 => x"53517288",
   273 => x"1381b72d",
   274 => x"8c127184",
   275 => x"2c708706",
   276 => x"55525272",
   277 => x"881381b7",
   278 => x"2d8c1271",
   279 => x"842c7087",
   280 => x"06555252",
   281 => x"72881381",
   282 => x"b72d7084",
   283 => x"2c708706",
   284 => x"51517094",
   285 => x"1381b72d",
   286 => x"028c050d",
   287 => x"0402d405",
   288 => x"0d7cb1d8",
   289 => x"525585f3",
   290 => x"2d9dc12d",
   291 => x"b7f80880",
   292 => x"2e83ae38",
   293 => x"86b52db7",
   294 => x"f8085390",
   295 => x"8a2db7f8",
   296 => x"0854b7f8",
   297 => x"08802e83",
   298 => x"9a38a1c4",
   299 => x"2db7f808",
   300 => x"802e8738",
   301 => x"b1f05189",
   302 => x"c70499ad",
   303 => x"2db7f808",
   304 => x"802ea238",
   305 => x"b2845185",
   306 => x"f32db29c",
   307 => x"5185f32d",
   308 => x"86942d72",
   309 => x"84075381",
   310 => x"0bfec40c",
   311 => x"72fec00c",
   312 => x"72518797",
   313 => x"2d840bfe",
   314 => x"c40cb2b8",
   315 => x"52b89851",
   316 => x"969c2d74",
   317 => x"822e0981",
   318 => x"06b738b7",
   319 => x"f808802e",
   320 => x"80e53872",
   321 => x"b8a40c87",
   322 => x"f62db7f8",
   323 => x"08b8a80c",
   324 => x"b8ac5480",
   325 => x"fd538074",
   326 => x"70840556",
   327 => x"0cff1353",
   328 => x"728025f2",
   329 => x"38b8a452",
   330 => x"b8985199",
   331 => x"872d8ae7",
   332 => x"0474812e",
   333 => x"098106af",
   334 => x"38b7f808",
   335 => x"802ea138",
   336 => x"b8a452b8",
   337 => x"985198e1",
   338 => x"2db8a408",
   339 => x"b8a80852",
   340 => x"5388b52d",
   341 => x"72fec00c",
   342 => x"72518797",
   343 => x"2d8ae704",
   344 => x"81eef751",
   345 => x"88b52db2",
   346 => x"c45185f3",
   347 => x"2db2dc52",
   348 => x"b8985196",
   349 => x"9c2db7f8",
   350 => x"089838b2",
   351 => x"e85185f3",
   352 => x"2db38052",
   353 => x"b8985196",
   354 => x"9c2db7f8",
   355 => x"08802e81",
   356 => x"b038b38c",
   357 => x"5185f32d",
   358 => x"b89c0857",
   359 => x"8077595a",
   360 => x"767a2e8b",
   361 => x"38811a78",
   362 => x"812a595a",
   363 => x"77f738f7",
   364 => x"1a5a8077",
   365 => x"25818038",
   366 => x"79527751",
   367 => x"84802db8",
   368 => x"a452b898",
   369 => x"5198e12d",
   370 => x"b7f80853",
   371 => x"b7f80880",
   372 => x"2e80c938",
   373 => x"b8a45b80",
   374 => x"598c8904",
   375 => x"7a708405",
   376 => x"5c087081",
   377 => x"ff067188",
   378 => x"2c7081ff",
   379 => x"0673902c",
   380 => x"7081ff06",
   381 => x"75982afe",
   382 => x"c80cfec8",
   383 => x"0c58fec8",
   384 => x"0c57fec8",
   385 => x"0c841a5a",
   386 => x"53765384",
   387 => x"80772584",
   388 => x"38848053",
   389 => x"727924c4",
   390 => x"388ca704",
   391 => x"b39c5185",
   392 => x"f32d7254",
   393 => x"8cc304b8",
   394 => x"985198b4",
   395 => x"2dfc8017",
   396 => x"81195957",
   397 => x"8bb20482",
   398 => x"0bfec40c",
   399 => x"81548cc3",
   400 => x"04805473",
   401 => x"b7f80c02",
   402 => x"ac050d04",
   403 => x"02f8050d",
   404 => x"a8972d81",
   405 => x"f72d8151",
   406 => x"84e52dfe",
   407 => x"c4528172",
   408 => x"0ca5902d",
   409 => x"a5902d84",
   410 => x"720c7351",
   411 => x"88fd2db4",
   412 => x"dc51a9f5",
   413 => x"2d805184",
   414 => x"e52d0288",
   415 => x"050d0402",
   416 => x"fc050d82",
   417 => x"518ccc2d",
   418 => x"0284050d",
   419 => x"0402fc05",
   420 => x"0d80518c",
   421 => x"cc2d0284",
   422 => x"050d0402",
   423 => x"ec050d84",
   424 => x"b8518797",
   425 => x"2d810bfe",
   426 => x"c40c84b8",
   427 => x"0bfec00c",
   428 => x"840bfec4",
   429 => x"0c830bfe",
   430 => x"cc0ca5ab",
   431 => x"2da88b2d",
   432 => x"a5902da5",
   433 => x"902d81f7",
   434 => x"2d815184",
   435 => x"e52da590",
   436 => x"2da5902d",
   437 => x"815184e5",
   438 => x"2d815188",
   439 => x"fd2db7f8",
   440 => x"08802e81",
   441 => x"d2388051",
   442 => x"84e52db4",
   443 => x"dc51a9f5",
   444 => x"2dbd8008",
   445 => x"8938bd84",
   446 => x"08802e80",
   447 => x"e238fed0",
   448 => x"08708106",
   449 => x"51527180",
   450 => x"2e80d438",
   451 => x"a8912dbd",
   452 => x"800870bd",
   453 => x"84087057",
   454 => x"55565280",
   455 => x"ff722584",
   456 => x"3880ff52",
   457 => x"80ff7325",
   458 => x"843880ff",
   459 => x"5371ff80",
   460 => x"258438ff",
   461 => x"805272ff",
   462 => x"80258438",
   463 => x"ff805374",
   464 => x"7231bd80",
   465 => x"0c737331",
   466 => x"bd840ca8",
   467 => x"8b2d7188",
   468 => x"2b83fe80",
   469 => x"067381ff",
   470 => x"067107fe",
   471 => x"d00c52a6",
   472 => x"902daa85",
   473 => x"2db7f808",
   474 => x"5386b52d",
   475 => x"b7f808fe",
   476 => x"c00c87f6",
   477 => x"2db7f808",
   478 => x"fed40c86",
   479 => x"b52db7f8",
   480 => x"08b89408",
   481 => x"2e9c38b7",
   482 => x"f808b894",
   483 => x"0c845272",
   484 => x"5184e52d",
   485 => x"a5902da5",
   486 => x"902dff12",
   487 => x"52718025",
   488 => x"ee387280",
   489 => x"2e89388a",
   490 => x"0bfec40c",
   491 => x"8df10482",
   492 => x"0bfec40c",
   493 => x"8df104b3",
   494 => x"ac5185f3",
   495 => x"2d820bfe",
   496 => x"c40c800b",
   497 => x"b7f80c02",
   498 => x"94050d04",
   499 => x"02e8050d",
   500 => x"77797b58",
   501 => x"55558053",
   502 => x"727625a3",
   503 => x"38747081",
   504 => x"055680f5",
   505 => x"2d747081",
   506 => x"055680f5",
   507 => x"2d525271",
   508 => x"712e8638",
   509 => x"81519081",
   510 => x"04811353",
   511 => x"8fd80480",
   512 => x"5170b7f8",
   513 => x"0c029805",
   514 => x"0d0402d8",
   515 => x"050d800b",
   516 => x"bcac0cb8",
   517 => x"a4528051",
   518 => x"a0a92db7",
   519 => x"f80854b7",
   520 => x"f8088c38",
   521 => x"b3c45185",
   522 => x"f32d7355",
   523 => x"95a50480",
   524 => x"56810bbc",
   525 => x"d00c8853",
   526 => x"b3d052b8",
   527 => x"da518fcc",
   528 => x"2db7f808",
   529 => x"762e0981",
   530 => x"068738b7",
   531 => x"f808bcd0",
   532 => x"0c8853b3",
   533 => x"dc52b8f6",
   534 => x"518fcc2d",
   535 => x"b7f80887",
   536 => x"38b7f808",
   537 => x"bcd00cbc",
   538 => x"d008802e",
   539 => x"80f638bb",
   540 => x"ea0b80f5",
   541 => x"2dbbeb0b",
   542 => x"80f52d71",
   543 => x"982b7190",
   544 => x"2b07bbec",
   545 => x"0b80f52d",
   546 => x"70882b72",
   547 => x"07bbed0b",
   548 => x"80f52d71",
   549 => x"07bca20b",
   550 => x"80f52dbc",
   551 => x"a30b80f5",
   552 => x"2d71882b",
   553 => x"07535f54",
   554 => x"525a5657",
   555 => x"557381ab",
   556 => x"aa2e0981",
   557 => x"068d3875",
   558 => x"51a1cb2d",
   559 => x"b7f80856",
   560 => x"91d00473",
   561 => x"82d4d52e",
   562 => x"8738b3e8",
   563 => x"51929104",
   564 => x"b8a45275",
   565 => x"51a0a92d",
   566 => x"b7f80855",
   567 => x"b7f80880",
   568 => x"2e83c238",
   569 => x"8853b3dc",
   570 => x"52b8f651",
   571 => x"8fcc2db7",
   572 => x"f8088938",
   573 => x"810bbcac",
   574 => x"0c929704",
   575 => x"8853b3d0",
   576 => x"52b8da51",
   577 => x"8fcc2db7",
   578 => x"f808802e",
   579 => x"8a38b3fc",
   580 => x"5185f32d",
   581 => x"92f104bc",
   582 => x"a20b80f5",
   583 => x"2d547380",
   584 => x"d52e0981",
   585 => x"0680ca38",
   586 => x"bca30b80",
   587 => x"f52d5473",
   588 => x"81aa2e09",
   589 => x"8106ba38",
   590 => x"800bb8a4",
   591 => x"0b80f52d",
   592 => x"56547481",
   593 => x"e92e8338",
   594 => x"81547481",
   595 => x"eb2e8c38",
   596 => x"80557375",
   597 => x"2e098106",
   598 => x"82cb38b8",
   599 => x"af0b80f5",
   600 => x"2d55748d",
   601 => x"38b8b00b",
   602 => x"80f52d54",
   603 => x"73822e86",
   604 => x"38805595",
   605 => x"a504b8b1",
   606 => x"0b80f52d",
   607 => x"70bca40c",
   608 => x"ff05bca8",
   609 => x"0cb8b20b",
   610 => x"80f52db8",
   611 => x"b30b80f5",
   612 => x"2d587605",
   613 => x"77828029",
   614 => x"0570bcb0",
   615 => x"0cb8b40b",
   616 => x"80f52d70",
   617 => x"bcc40cbc",
   618 => x"ac085957",
   619 => x"5876802e",
   620 => x"81a33888",
   621 => x"53b3dc52",
   622 => x"b8f6518f",
   623 => x"cc2db7f8",
   624 => x"0881e238",
   625 => x"bca40870",
   626 => x"842bbcc8",
   627 => x"0c70bcc0",
   628 => x"0cb8c90b",
   629 => x"80f52db8",
   630 => x"c80b80f5",
   631 => x"2d718280",
   632 => x"2905b8ca",
   633 => x"0b80f52d",
   634 => x"70848080",
   635 => x"2912b8cb",
   636 => x"0b80f52d",
   637 => x"7081800a",
   638 => x"291270bc",
   639 => x"cc0cbcc4",
   640 => x"087129bc",
   641 => x"b0080570",
   642 => x"bcb40cb8",
   643 => x"d10b80f5",
   644 => x"2db8d00b",
   645 => x"80f52d71",
   646 => x"82802905",
   647 => x"b8d20b80",
   648 => x"f52d7084",
   649 => x"80802912",
   650 => x"b8d30b80",
   651 => x"f52d7098",
   652 => x"2b81f00a",
   653 => x"06720570",
   654 => x"bcb80cfe",
   655 => x"117e2977",
   656 => x"05bcbc0c",
   657 => x"52595243",
   658 => x"545e5152",
   659 => x"59525d57",
   660 => x"595795a3",
   661 => x"04b8b60b",
   662 => x"80f52db8",
   663 => x"b50b80f5",
   664 => x"2d718280",
   665 => x"290570bc",
   666 => x"c80c70a0",
   667 => x"2983ff05",
   668 => x"70892a70",
   669 => x"bcc00cb8",
   670 => x"bb0b80f5",
   671 => x"2db8ba0b",
   672 => x"80f52d71",
   673 => x"82802905",
   674 => x"70bccc0c",
   675 => x"7b71291e",
   676 => x"70bcbc0c",
   677 => x"7dbcb80c",
   678 => x"7305bcb4",
   679 => x"0c555e51",
   680 => x"51555581",
   681 => x"5574b7f8",
   682 => x"0c02a805",
   683 => x"0d0402ec",
   684 => x"050d7670",
   685 => x"872c7180",
   686 => x"ff065556",
   687 => x"54bcac08",
   688 => x"8a387388",
   689 => x"2c7481ff",
   690 => x"065455b8",
   691 => x"a452bcb0",
   692 => x"081551a0",
   693 => x"a92db7f8",
   694 => x"0854b7f8",
   695 => x"08802eb3",
   696 => x"38bcac08",
   697 => x"802e9838",
   698 => x"728429b8",
   699 => x"a4057008",
   700 => x"5253a1cb",
   701 => x"2db7f808",
   702 => x"f00a0653",
   703 => x"96910472",
   704 => x"10b8a405",
   705 => x"7080e02d",
   706 => x"5253a1fb",
   707 => x"2db7f808",
   708 => x"53725473",
   709 => x"b7f80c02",
   710 => x"94050d04",
   711 => x"02c8050d",
   712 => x"7f615f5b",
   713 => x"800bbcb8",
   714 => x"08bcbc08",
   715 => x"595d56bc",
   716 => x"ac08762e",
   717 => x"8a38bca4",
   718 => x"08842b58",
   719 => x"96c504bc",
   720 => x"c008842b",
   721 => x"58805978",
   722 => x"782781a9",
   723 => x"38788f06",
   724 => x"a0175754",
   725 => x"738f38b8",
   726 => x"a4527651",
   727 => x"811757a0",
   728 => x"a92db8a4",
   729 => x"56807680",
   730 => x"f52d5654",
   731 => x"74742e83",
   732 => x"38815474",
   733 => x"81e52e80",
   734 => x"f6388170",
   735 => x"7506555d",
   736 => x"73802e80",
   737 => x"ea388b16",
   738 => x"80f52d98",
   739 => x"065a7980",
   740 => x"de388b53",
   741 => x"7d527551",
   742 => x"8fcc2db7",
   743 => x"f80880cf",
   744 => x"389c1608",
   745 => x"51a1cb2d",
   746 => x"b7f80884",
   747 => x"1c0c9a16",
   748 => x"80e02d51",
   749 => x"a1fb2db7",
   750 => x"f808b7f8",
   751 => x"08881d0c",
   752 => x"b7f80855",
   753 => x"55bcac08",
   754 => x"802e9838",
   755 => x"941680e0",
   756 => x"2d51a1fb",
   757 => x"2db7f808",
   758 => x"902b83ff",
   759 => x"f00a0670",
   760 => x"16515473",
   761 => x"881c0c79",
   762 => x"7b0c7c54",
   763 => x"98ab0481",
   764 => x"195996c7",
   765 => x"04bcac08",
   766 => x"802eae38",
   767 => x"7b5195ae",
   768 => x"2db7f808",
   769 => x"b7f80880",
   770 => x"fffffff8",
   771 => x"06555c73",
   772 => x"80ffffff",
   773 => x"f82e9238",
   774 => x"b7f808fe",
   775 => x"05bca408",
   776 => x"29bcb408",
   777 => x"055796c5",
   778 => x"04805473",
   779 => x"b7f80c02",
   780 => x"b8050d04",
   781 => x"02f4050d",
   782 => x"74700881",
   783 => x"05710c70",
   784 => x"08bca808",
   785 => x"06535371",
   786 => x"8e388813",
   787 => x"085195ae",
   788 => x"2db7f808",
   789 => x"88140c81",
   790 => x"0bb7f80c",
   791 => x"028c050d",
   792 => x"0402f005",
   793 => x"0d758811",
   794 => x"08fe05bc",
   795 => x"a40829bc",
   796 => x"b4081172",
   797 => x"08bca808",
   798 => x"06057955",
   799 => x"535454a0",
   800 => x"a92d0290",
   801 => x"050d0402",
   802 => x"f0050d75",
   803 => x"881108fe",
   804 => x"05bca408",
   805 => x"29bcb408",
   806 => x"117208bc",
   807 => x"a8080605",
   808 => x"79555354",
   809 => x"549ee92d",
   810 => x"0290050d",
   811 => x"04bcac08",
   812 => x"b7f80c04",
   813 => x"02f4050d",
   814 => x"d45281ff",
   815 => x"720c7108",
   816 => x"5381ff72",
   817 => x"0c72882b",
   818 => x"83fe8006",
   819 => x"72087081",
   820 => x"ff065152",
   821 => x"5381ff72",
   822 => x"0c727107",
   823 => x"882b7208",
   824 => x"7081ff06",
   825 => x"51525381",
   826 => x"ff720c72",
   827 => x"7107882b",
   828 => x"72087081",
   829 => x"ff067207",
   830 => x"b7f80c52",
   831 => x"53028c05",
   832 => x"0d0402f4",
   833 => x"050d7476",
   834 => x"7181ff06",
   835 => x"d40c5353",
   836 => x"bcd40885",
   837 => x"3871892b",
   838 => x"5271982a",
   839 => x"d40c7190",
   840 => x"2a7081ff",
   841 => x"06d40c51",
   842 => x"71882a70",
   843 => x"81ff06d4",
   844 => x"0c517181",
   845 => x"ff06d40c",
   846 => x"72902a70",
   847 => x"81ff06d4",
   848 => x"0c51d408",
   849 => x"7081ff06",
   850 => x"515182b8",
   851 => x"bf527081",
   852 => x"ff2e0981",
   853 => x"06943881",
   854 => x"ff0bd40c",
   855 => x"d4087081",
   856 => x"ff06ff14",
   857 => x"54515171",
   858 => x"e53870b7",
   859 => x"f80c028c",
   860 => x"050d0402",
   861 => x"fc050d81",
   862 => x"c75181ff",
   863 => x"0bd40cff",
   864 => x"11517080",
   865 => x"25f43802",
   866 => x"84050d04",
   867 => x"02f0050d",
   868 => x"9af32d8f",
   869 => x"cf538052",
   870 => x"87fc80f7",
   871 => x"519a822d",
   872 => x"b7f80854",
   873 => x"b7f80881",
   874 => x"2e098106",
   875 => x"a33881ff",
   876 => x"0bd40c82",
   877 => x"0a52849c",
   878 => x"80e9519a",
   879 => x"822db7f8",
   880 => x"088b3881",
   881 => x"ff0bd40c",
   882 => x"73539bd6",
   883 => x"049af32d",
   884 => x"ff135372",
   885 => x"c13872b7",
   886 => x"f80c0290",
   887 => x"050d0402",
   888 => x"f4050d81",
   889 => x"ff0bd40c",
   890 => x"93538052",
   891 => x"87fc80c1",
   892 => x"519a822d",
   893 => x"b7f8088b",
   894 => x"3881ff0b",
   895 => x"d40c8153",
   896 => x"9c8c049a",
   897 => x"f32dff13",
   898 => x"5372df38",
   899 => x"72b7f80c",
   900 => x"028c050d",
   901 => x"0402f005",
   902 => x"0d9af32d",
   903 => x"83aa5284",
   904 => x"9c80c851",
   905 => x"9a822db7",
   906 => x"f808812e",
   907 => x"09810692",
   908 => x"3899b42d",
   909 => x"b7f80883",
   910 => x"ffff0653",
   911 => x"7283aa2e",
   912 => x"97389bdf",
   913 => x"2d9cd304",
   914 => x"81549db8",
   915 => x"04b48851",
   916 => x"85f32d80",
   917 => x"549db804",
   918 => x"81ff0bd4",
   919 => x"0cb1539b",
   920 => x"8c2db7f8",
   921 => x"08802e80",
   922 => x"c0388052",
   923 => x"87fc80fa",
   924 => x"519a822d",
   925 => x"b7f808b1",
   926 => x"3881ff0b",
   927 => x"d40cd408",
   928 => x"5381ff0b",
   929 => x"d40c81ff",
   930 => x"0bd40c81",
   931 => x"ff0bd40c",
   932 => x"81ff0bd4",
   933 => x"0c72862a",
   934 => x"708106b7",
   935 => x"f8085651",
   936 => x"5372802e",
   937 => x"93389cc8",
   938 => x"0472822e",
   939 => x"ff9f38ff",
   940 => x"135372ff",
   941 => x"aa387254",
   942 => x"73b7f80c",
   943 => x"0290050d",
   944 => x"0402f005",
   945 => x"0d810bbc",
   946 => x"d40c8454",
   947 => x"d008708f",
   948 => x"2a708106",
   949 => x"51515372",
   950 => x"f33872d0",
   951 => x"0c9af32d",
   952 => x"b4985185",
   953 => x"f32dd008",
   954 => x"708f2a70",
   955 => x"81065151",
   956 => x"5372f338",
   957 => x"810bd00c",
   958 => x"b1538052",
   959 => x"84d480c0",
   960 => x"519a822d",
   961 => x"b7f80881",
   962 => x"2ea13872",
   963 => x"822e0981",
   964 => x"068c38b4",
   965 => x"a45185f3",
   966 => x"2d80539e",
   967 => x"e004ff13",
   968 => x"5372d738",
   969 => x"ff145473",
   970 => x"ffa2389c",
   971 => x"952db7f8",
   972 => x"08bcd40c",
   973 => x"b7f8088b",
   974 => x"38815287",
   975 => x"fc80d051",
   976 => x"9a822d81",
   977 => x"ff0bd40c",
   978 => x"d008708f",
   979 => x"2a708106",
   980 => x"51515372",
   981 => x"f33872d0",
   982 => x"0c81ff0b",
   983 => x"d40c8153",
   984 => x"72b7f80c",
   985 => x"0290050d",
   986 => x"0402e805",
   987 => x"0d785681",
   988 => x"ff0bd40c",
   989 => x"d008708f",
   990 => x"2a708106",
   991 => x"51515372",
   992 => x"f3388281",
   993 => x"0bd00c81",
   994 => x"ff0bd40c",
   995 => x"775287fc",
   996 => x"80d8519a",
   997 => x"822db7f8",
   998 => x"08802e8c",
   999 => x"38b4bc51",
  1000 => x"85f32d81",
  1001 => x"53a0a004",
  1002 => x"81ff0bd4",
  1003 => x"0c81fe0b",
  1004 => x"d40c80ff",
  1005 => x"55757084",
  1006 => x"05570870",
  1007 => x"982ad40c",
  1008 => x"70902c70",
  1009 => x"81ff06d4",
  1010 => x"0c547088",
  1011 => x"2c7081ff",
  1012 => x"06d40c54",
  1013 => x"7081ff06",
  1014 => x"d40c54ff",
  1015 => x"15557480",
  1016 => x"25d33881",
  1017 => x"ff0bd40c",
  1018 => x"81ff0bd4",
  1019 => x"0c81ff0b",
  1020 => x"d40c868d",
  1021 => x"a05481ff",
  1022 => x"0bd40cd4",
  1023 => x"0881ff06",
  1024 => x"55748738",
  1025 => x"ff145473",
  1026 => x"ed3881ff",
  1027 => x"0bd40cd0",
  1028 => x"08708f2a",
  1029 => x"70810651",
  1030 => x"515372f3",
  1031 => x"3872d00c",
  1032 => x"72b7f80c",
  1033 => x"0298050d",
  1034 => x"0402e805",
  1035 => x"0d785580",
  1036 => x"5681ff0b",
  1037 => x"d40cd008",
  1038 => x"708f2a70",
  1039 => x"81065151",
  1040 => x"5372f338",
  1041 => x"82810bd0",
  1042 => x"0c81ff0b",
  1043 => x"d40c7752",
  1044 => x"87fc80d1",
  1045 => x"519a822d",
  1046 => x"80dbc6df",
  1047 => x"54b7f808",
  1048 => x"802e8a38",
  1049 => x"b39c5185",
  1050 => x"f32da1bb",
  1051 => x"0481ff0b",
  1052 => x"d40cd408",
  1053 => x"7081ff06",
  1054 => x"51537281",
  1055 => x"fe2e0981",
  1056 => x"069d3880",
  1057 => x"ff5399b4",
  1058 => x"2db7f808",
  1059 => x"75708405",
  1060 => x"570cff13",
  1061 => x"53728025",
  1062 => x"ed388156",
  1063 => x"a1a504ff",
  1064 => x"145473c9",
  1065 => x"3881ff0b",
  1066 => x"d40cd008",
  1067 => x"708f2a70",
  1068 => x"81065151",
  1069 => x"5372f338",
  1070 => x"72d00c75",
  1071 => x"b7f80c02",
  1072 => x"98050d04",
  1073 => x"bcd408b7",
  1074 => x"f80c0402",
  1075 => x"f4050d74",
  1076 => x"70882a83",
  1077 => x"fe800670",
  1078 => x"72982a07",
  1079 => x"72882b87",
  1080 => x"fc808006",
  1081 => x"73982b81",
  1082 => x"f00a0671",
  1083 => x"730707b7",
  1084 => x"f80c5651",
  1085 => x"5351028c",
  1086 => x"050d0402",
  1087 => x"f8050d02",
  1088 => x"8e0580f5",
  1089 => x"2d74882b",
  1090 => x"077083ff",
  1091 => x"ff06b7f8",
  1092 => x"0c510288",
  1093 => x"050d0402",
  1094 => x"fc050d72",
  1095 => x"5180710c",
  1096 => x"800b8412",
  1097 => x"0c028405",
  1098 => x"0d0402f0",
  1099 => x"050d7570",
  1100 => x"08841208",
  1101 => x"535353ff",
  1102 => x"5471712e",
  1103 => x"a838a891",
  1104 => x"2d841308",
  1105 => x"70842914",
  1106 => x"88117008",
  1107 => x"7081ff06",
  1108 => x"84180881",
  1109 => x"11870684",
  1110 => x"1a0c5351",
  1111 => x"55515151",
  1112 => x"a88b2d71",
  1113 => x"5473b7f8",
  1114 => x"0c029005",
  1115 => x"0d0402f4",
  1116 => x"050da891",
  1117 => x"2de008e4",
  1118 => x"08718b2a",
  1119 => x"70810651",
  1120 => x"53545270",
  1121 => x"802e9d38",
  1122 => x"bcd80870",
  1123 => x"8429bce0",
  1124 => x"057381ff",
  1125 => x"06710c51",
  1126 => x"51bcd808",
  1127 => x"81118706",
  1128 => x"bcd80c51",
  1129 => x"728b2a70",
  1130 => x"81065151",
  1131 => x"70802e81",
  1132 => x"9238b7a8",
  1133 => x"088429bd",
  1134 => x"8c057381",
  1135 => x"ff06710c",
  1136 => x"51b7a808",
  1137 => x"8105b7a8",
  1138 => x"0c850bb7",
  1139 => x"a40cb7a8",
  1140 => x"08b7a008",
  1141 => x"2e098106",
  1142 => x"81a63880",
  1143 => x"0bb7a80c",
  1144 => x"bd9c0881",
  1145 => x"9b38bd8c",
  1146 => x"08700970",
  1147 => x"8306fecc",
  1148 => x"0c527085",
  1149 => x"2a708106",
  1150 => x"bd840855",
  1151 => x"51525370",
  1152 => x"802e8e38",
  1153 => x"bd9408fe",
  1154 => x"803212bd",
  1155 => x"840ca498",
  1156 => x"04bd9408",
  1157 => x"12bd840c",
  1158 => x"72842a70",
  1159 => x"8106bd80",
  1160 => x"08545151",
  1161 => x"70802e90",
  1162 => x"38bd9008",
  1163 => x"81ff3212",
  1164 => x"8105bd80",
  1165 => x"0ca58004",
  1166 => x"71bd9008",
  1167 => x"31bd800c",
  1168 => x"a58004b7",
  1169 => x"a408ff05",
  1170 => x"b7a40cb7",
  1171 => x"a408ff2e",
  1172 => x"098106ac",
  1173 => x"38b7a808",
  1174 => x"802e9238",
  1175 => x"810bbd9c",
  1176 => x"0c870bb7",
  1177 => x"a00831b7",
  1178 => x"a00ca4fb",
  1179 => x"04bd9c08",
  1180 => x"5170802e",
  1181 => x"8638ff11",
  1182 => x"bd9c0c80",
  1183 => x"0bb7a80c",
  1184 => x"800bbd88",
  1185 => x"0ca8842d",
  1186 => x"a88b2d02",
  1187 => x"8c050d04",
  1188 => x"02fc050d",
  1189 => x"a8912d81",
  1190 => x"0bbd880c",
  1191 => x"a88b2dbd",
  1192 => x"88085170",
  1193 => x"fa380284",
  1194 => x"050d0402",
  1195 => x"f8050dbc",
  1196 => x"d851a297",
  1197 => x"2d800bbd",
  1198 => x"9c0c830b",
  1199 => x"b7a00ce4",
  1200 => x"08708c2a",
  1201 => x"70810651",
  1202 => x"51527180",
  1203 => x"2e863884",
  1204 => x"0bb7a00c",
  1205 => x"e408708d",
  1206 => x"2a708106",
  1207 => x"51515271",
  1208 => x"802e9f38",
  1209 => x"870bb7a0",
  1210 => x"0831b7a0",
  1211 => x"0ce40870",
  1212 => x"8a2a7081",
  1213 => x"06515152",
  1214 => x"71802ef1",
  1215 => x"3881f40b",
  1216 => x"e40ca2ee",
  1217 => x"51a8802d",
  1218 => x"a7aa2d02",
  1219 => x"88050d04",
  1220 => x"02f4050d",
  1221 => x"a79204b7",
  1222 => x"f80881f0",
  1223 => x"2e098106",
  1224 => x"8938810b",
  1225 => x"b7ec0ca7",
  1226 => x"9204b7f8",
  1227 => x"0881e02e",
  1228 => x"09810689",
  1229 => x"38810bb7",
  1230 => x"f00ca792",
  1231 => x"04b7f808",
  1232 => x"52b7f008",
  1233 => x"802e8838",
  1234 => x"b7f80881",
  1235 => x"80055271",
  1236 => x"842c728f",
  1237 => x"065353b7",
  1238 => x"ec08802e",
  1239 => x"99387284",
  1240 => x"29b7ac05",
  1241 => x"72138171",
  1242 => x"2b700973",
  1243 => x"0806730c",
  1244 => x"515353a7",
  1245 => x"88047284",
  1246 => x"29b7ac05",
  1247 => x"72138371",
  1248 => x"2b720807",
  1249 => x"720c5353",
  1250 => x"800bb7f0",
  1251 => x"0c800bb7",
  1252 => x"ec0cbcd8",
  1253 => x"51a2aa2d",
  1254 => x"b7f808ff",
  1255 => x"24fef838",
  1256 => x"800bb7f8",
  1257 => x"0c028c05",
  1258 => x"0d0402f8",
  1259 => x"050db7ac",
  1260 => x"528f5180",
  1261 => x"72708405",
  1262 => x"540cff11",
  1263 => x"51708025",
  1264 => x"f2380288",
  1265 => x"050d0402",
  1266 => x"f0050d75",
  1267 => x"51a8912d",
  1268 => x"70822cfc",
  1269 => x"06b7ac11",
  1270 => x"72109e06",
  1271 => x"71087072",
  1272 => x"2a708306",
  1273 => x"82742b70",
  1274 => x"09740676",
  1275 => x"0c545156",
  1276 => x"57535153",
  1277 => x"a88b2d71",
  1278 => x"b7f80c02",
  1279 => x"90050d04",
  1280 => x"71980c04",
  1281 => x"ffb008b7",
  1282 => x"f80c0481",
  1283 => x"0bffb00c",
  1284 => x"04800bff",
  1285 => x"b00c0402",
  1286 => x"fc050d80",
  1287 => x"0bb7f40c",
  1288 => x"805184e5",
  1289 => x"2d028405",
  1290 => x"0d0402ec",
  1291 => x"050d7654",
  1292 => x"8052870b",
  1293 => x"881580f5",
  1294 => x"2d565374",
  1295 => x"72248338",
  1296 => x"a0537251",
  1297 => x"82ee2d81",
  1298 => x"128b1580",
  1299 => x"f52d5452",
  1300 => x"727225de",
  1301 => x"38029405",
  1302 => x"0d0402f0",
  1303 => x"050dbda4",
  1304 => x"085481f7",
  1305 => x"2d800bbd",
  1306 => x"a80c7308",
  1307 => x"802e8180",
  1308 => x"38820bb8",
  1309 => x"8c0cbda8",
  1310 => x"088f06b8",
  1311 => x"880c7308",
  1312 => x"5271832e",
  1313 => x"96387183",
  1314 => x"26893871",
  1315 => x"812eaf38",
  1316 => x"a9db0471",
  1317 => x"852e9f38",
  1318 => x"a9db0488",
  1319 => x"1480f52d",
  1320 => x"841508b4",
  1321 => x"cc535452",
  1322 => x"85f32d71",
  1323 => x"84291370",
  1324 => x"085252a9",
  1325 => x"df047351",
  1326 => x"a8aa2da9",
  1327 => x"db04bda0",
  1328 => x"08881508",
  1329 => x"2c708106",
  1330 => x"51527180",
  1331 => x"2e8738b4",
  1332 => x"d051a9d8",
  1333 => x"04b4d451",
  1334 => x"85f32d84",
  1335 => x"14085185",
  1336 => x"f32dbda8",
  1337 => x"088105bd",
  1338 => x"a80c8c14",
  1339 => x"54a8ea04",
  1340 => x"0290050d",
  1341 => x"0471bda4",
  1342 => x"0ca8da2d",
  1343 => x"bda808ff",
  1344 => x"05bdac0c",
  1345 => x"0402ec05",
  1346 => x"0dbda408",
  1347 => x"5580f851",
  1348 => x"a7c72db7",
  1349 => x"f808812a",
  1350 => x"70810651",
  1351 => x"52719b38",
  1352 => x"8751a7c7",
  1353 => x"2db7f808",
  1354 => x"812a7081",
  1355 => x"06515271",
  1356 => x"802eb138",
  1357 => x"aaba04a6",
  1358 => x"902d8751",
  1359 => x"a7c72db7",
  1360 => x"f808f438",
  1361 => x"aaca04a6",
  1362 => x"902d80f8",
  1363 => x"51a7c72d",
  1364 => x"b7f808f3",
  1365 => x"38b7f408",
  1366 => x"813270b7",
  1367 => x"f40c7052",
  1368 => x"5284e52d",
  1369 => x"b7f408a2",
  1370 => x"3880da51",
  1371 => x"a7c72d81",
  1372 => x"f551a7c7",
  1373 => x"2d81f251",
  1374 => x"a7c72d81",
  1375 => x"eb51a7c7",
  1376 => x"2d81f451",
  1377 => x"a7c72dae",
  1378 => x"ce0481f5",
  1379 => x"51a7c72d",
  1380 => x"b7f80881",
  1381 => x"2a708106",
  1382 => x"51527180",
  1383 => x"2e8f38bd",
  1384 => x"ac085271",
  1385 => x"802e8638",
  1386 => x"ff12bdac",
  1387 => x"0c81f251",
  1388 => x"a7c72db7",
  1389 => x"f808812a",
  1390 => x"70810651",
  1391 => x"5271802e",
  1392 => x"9538bda8",
  1393 => x"08ff05bd",
  1394 => x"ac085452",
  1395 => x"72722586",
  1396 => x"388113bd",
  1397 => x"ac0cbdac",
  1398 => x"08705354",
  1399 => x"73802e8a",
  1400 => x"388c15ff",
  1401 => x"155555ab",
  1402 => x"dc04820b",
  1403 => x"b88c0c71",
  1404 => x"8f06b888",
  1405 => x"0c81eb51",
  1406 => x"a7c72db7",
  1407 => x"f808812a",
  1408 => x"70810651",
  1409 => x"5271802e",
  1410 => x"ad387408",
  1411 => x"852e0981",
  1412 => x"06a43888",
  1413 => x"1580f52d",
  1414 => x"ff055271",
  1415 => x"881681b7",
  1416 => x"2d71982b",
  1417 => x"52718025",
  1418 => x"8838800b",
  1419 => x"881681b7",
  1420 => x"2d7451a8",
  1421 => x"aa2d81f4",
  1422 => x"51a7c72d",
  1423 => x"b7f80881",
  1424 => x"2a708106",
  1425 => x"51527180",
  1426 => x"2eb33874",
  1427 => x"08852e09",
  1428 => x"8106aa38",
  1429 => x"881580f5",
  1430 => x"2d810552",
  1431 => x"71881681",
  1432 => x"b72d7181",
  1433 => x"ff068b16",
  1434 => x"80f52d54",
  1435 => x"52727227",
  1436 => x"87387288",
  1437 => x"1681b72d",
  1438 => x"7451a8aa",
  1439 => x"2d80da51",
  1440 => x"a7c72db7",
  1441 => x"f808812a",
  1442 => x"70810651",
  1443 => x"5271802e",
  1444 => x"80fb38bd",
  1445 => x"a408bdac",
  1446 => x"08555373",
  1447 => x"802e8a38",
  1448 => x"8c13ff15",
  1449 => x"5553ad9b",
  1450 => x"04720852",
  1451 => x"71822ea6",
  1452 => x"38718226",
  1453 => x"89387181",
  1454 => x"2ea538ae",
  1455 => x"8d047183",
  1456 => x"2ead3871",
  1457 => x"842e0981",
  1458 => x"0680c238",
  1459 => x"88130851",
  1460 => x"a9f52dae",
  1461 => x"8d048813",
  1462 => x"0852712d",
  1463 => x"ae8d0481",
  1464 => x"0b881408",
  1465 => x"2bbda008",
  1466 => x"32bda00c",
  1467 => x"ae8a0488",
  1468 => x"1380f52d",
  1469 => x"81058b14",
  1470 => x"80f52d53",
  1471 => x"54717424",
  1472 => x"83388054",
  1473 => x"73881481",
  1474 => x"b72da8da",
  1475 => x"2d805480",
  1476 => x"0bb88c0c",
  1477 => x"738f06b8",
  1478 => x"880ca052",
  1479 => x"73bdac08",
  1480 => x"2e098106",
  1481 => x"9838bda8",
  1482 => x"08ff0574",
  1483 => x"32700981",
  1484 => x"05707207",
  1485 => x"9f2a9171",
  1486 => x"31515153",
  1487 => x"53715182",
  1488 => x"ee2d8114",
  1489 => x"548e7425",
  1490 => x"c638b7f4",
  1491 => x"085271b7",
  1492 => x"f80c0294",
  1493 => x"050d0400",
  1494 => x"00ffffff",
  1495 => x"ff00ffff",
  1496 => x"ffff00ff",
  1497 => x"ffffff00",
  1498 => x"52657365",
  1499 => x"74000000",
  1500 => x"53617665",
  1501 => x"20616e64",
  1502 => x"20526573",
  1503 => x"65740000",
  1504 => x"4f707469",
  1505 => x"6f6e7320",
  1506 => x"10000000",
  1507 => x"536f756e",
  1508 => x"64201000",
  1509 => x"54757262",
  1510 => x"6f000000",
  1511 => x"4d6f7573",
  1512 => x"6520656d",
  1513 => x"756c6174",
  1514 => x"696f6e00",
  1515 => x"45786974",
  1516 => x"00000000",
  1517 => x"4d617374",
  1518 => x"65720000",
  1519 => x"4f504c4c",
  1520 => x"00000000",
  1521 => x"53434300",
  1522 => x"50534700",
  1523 => x"4261636b",
  1524 => x"00000000",
  1525 => x"5363616e",
  1526 => x"6c696e65",
  1527 => x"73000000",
  1528 => x"53442043",
  1529 => x"61726400",
  1530 => x"4a617061",
  1531 => x"6e657365",
  1532 => x"206b6579",
  1533 => x"206c6179",
  1534 => x"6f757400",
  1535 => x"32303438",
  1536 => x"4b422052",
  1537 => x"414d0000",
  1538 => x"34303936",
  1539 => x"4b422052",
  1540 => x"414d0000",
  1541 => x"536c323a",
  1542 => x"204e6f6e",
  1543 => x"65000000",
  1544 => x"536c323a",
  1545 => x"20455345",
  1546 => x"2d534343",
  1547 => x"20314d42",
  1548 => x"2f534343",
  1549 => x"2d490000",
  1550 => x"536c323a",
  1551 => x"20455345",
  1552 => x"2d52414d",
  1553 => x"20314d42",
  1554 => x"2f415343",
  1555 => x"49493800",
  1556 => x"536c323a",
  1557 => x"20455345",
  1558 => x"2d52414d",
  1559 => x"20314d42",
  1560 => x"2f415343",
  1561 => x"49493136",
  1562 => x"00000000",
  1563 => x"536c313a",
  1564 => x"204e6f6e",
  1565 => x"65000000",
  1566 => x"536c313a",
  1567 => x"20455345",
  1568 => x"2d534343",
  1569 => x"20314d42",
  1570 => x"2f534343",
  1571 => x"2d490000",
  1572 => x"536c313a",
  1573 => x"204d6567",
  1574 => x"6152414d",
  1575 => x"00000000",
  1576 => x"56474120",
  1577 => x"2d203331",
  1578 => x"4b487a2c",
  1579 => x"20363048",
  1580 => x"7a000000",
  1581 => x"56474120",
  1582 => x"2d203331",
  1583 => x"4b487a2c",
  1584 => x"20353048",
  1585 => x"7a000000",
  1586 => x"5456202d",
  1587 => x"20343830",
  1588 => x"692c2036",
  1589 => x"30487a00",
  1590 => x"496e6974",
  1591 => x"69616c69",
  1592 => x"7a696e67",
  1593 => x"20534420",
  1594 => x"63617264",
  1595 => x"0a000000",
  1596 => x"53444843",
  1597 => x"206e6f74",
  1598 => x"20737570",
  1599 => x"706f7274",
  1600 => x"65643b00",
  1601 => x"46617433",
  1602 => x"32206e6f",
  1603 => x"74207375",
  1604 => x"70706f72",
  1605 => x"7465643b",
  1606 => x"00000000",
  1607 => x"0a646973",
  1608 => x"61626c69",
  1609 => x"6e672053",
  1610 => x"44206361",
  1611 => x"72640a10",
  1612 => x"204f4b0a",
  1613 => x"00000000",
  1614 => x"4f434d53",
  1615 => x"58202020",
  1616 => x"43464700",
  1617 => x"54727969",
  1618 => x"6e67204d",
  1619 => x"53583342",
  1620 => x"494f532e",
  1621 => x"5359530a",
  1622 => x"00000000",
  1623 => x"4d535833",
  1624 => x"42494f53",
  1625 => x"53595300",
  1626 => x"54727969",
  1627 => x"6e672042",
  1628 => x"494f535f",
  1629 => x"4d32502e",
  1630 => x"524f4d0a",
  1631 => x"00000000",
  1632 => x"42494f53",
  1633 => x"5f4d3250",
  1634 => x"524f4d00",
  1635 => x"4c6f6164",
  1636 => x"696e6720",
  1637 => x"42494f53",
  1638 => x"0a000000",
  1639 => x"52656164",
  1640 => x"20666169",
  1641 => x"6c65640a",
  1642 => x"00000000",
  1643 => x"4c6f6164",
  1644 => x"696e6720",
  1645 => x"42494f53",
  1646 => x"20666169",
  1647 => x"6c65640a",
  1648 => x"00000000",
  1649 => x"4d425220",
  1650 => x"6661696c",
  1651 => x"0a000000",
  1652 => x"46415431",
  1653 => x"36202020",
  1654 => x"00000000",
  1655 => x"46415433",
  1656 => x"32202020",
  1657 => x"00000000",
  1658 => x"4e6f2070",
  1659 => x"61727469",
  1660 => x"74696f6e",
  1661 => x"20736967",
  1662 => x"0a000000",
  1663 => x"42616420",
  1664 => x"70617274",
  1665 => x"0a000000",
  1666 => x"53444843",
  1667 => x"20657272",
  1668 => x"6f72210a",
  1669 => x"00000000",
  1670 => x"53442069",
  1671 => x"6e69742e",
  1672 => x"2e2e0a00",
  1673 => x"53442063",
  1674 => x"61726420",
  1675 => x"72657365",
  1676 => x"74206661",
  1677 => x"696c6564",
  1678 => x"210a0000",
  1679 => x"57726974",
  1680 => x"65206661",
  1681 => x"696c6564",
  1682 => x"0a000000",
  1683 => x"16200000",
  1684 => x"14200000",
  1685 => x"15200000",
  1686 => x"00000002",
  1687 => x"00000002",
  1688 => x"00001768",
  1689 => x"0000068d",
  1690 => x"00000002",
  1691 => x"00001770",
  1692 => x"0000067f",
  1693 => x"00000004",
  1694 => x"00001780",
  1695 => x"00001b04",
  1696 => x"00000004",
  1697 => x"0000178c",
  1698 => x"00001abc",
  1699 => x"00000001",
  1700 => x"00001794",
  1701 => x"00000007",
  1702 => x"00000001",
  1703 => x"0000179c",
  1704 => x"0000000a",
  1705 => x"00000002",
  1706 => x"000017ac",
  1707 => x"00001417",
  1708 => x"00000000",
  1709 => x"00000000",
  1710 => x"00000000",
  1711 => x"00000005",
  1712 => x"000017b4",
  1713 => x"00000007",
  1714 => x"00000005",
  1715 => x"000017bc",
  1716 => x"00000007",
  1717 => x"00000005",
  1718 => x"000017c4",
  1719 => x"00000007",
  1720 => x"00000005",
  1721 => x"000017c8",
  1722 => x"00000007",
  1723 => x"00000004",
  1724 => x"000017cc",
  1725 => x"00001a5c",
  1726 => x"00000000",
  1727 => x"00000000",
  1728 => x"00000000",
  1729 => x"00000003",
  1730 => x"00001b94",
  1731 => x"00000003",
  1732 => x"00000001",
  1733 => x"000017d4",
  1734 => x"0000000b",
  1735 => x"00000001",
  1736 => x"000017e0",
  1737 => x"00000002",
  1738 => x"00000003",
  1739 => x"00001b88",
  1740 => x"00000003",
  1741 => x"00000003",
  1742 => x"00001b78",
  1743 => x"00000004",
  1744 => x"00000001",
  1745 => x"000017e8",
  1746 => x"00000006",
  1747 => x"00000003",
  1748 => x"00001b70",
  1749 => x"00000002",
  1750 => x"00000004",
  1751 => x"000017cc",
  1752 => x"00001a5c",
  1753 => x"00000000",
  1754 => x"00000000",
  1755 => x"00000000",
  1756 => x"000017fc",
  1757 => x"00001808",
  1758 => x"00001814",
  1759 => x"00001820",
  1760 => x"00001838",
  1761 => x"00001850",
  1762 => x"0000186c",
  1763 => x"00001878",
  1764 => x"00001890",
  1765 => x"000018a0",
  1766 => x"000018b4",
  1767 => x"000018c8",
  1768 => x"00000003",
  1769 => x"00000000",
  1770 => x"00000000",
  1771 => x"00000000",
  1772 => x"00000000",
  1773 => x"00000000",
  1774 => x"00000000",
  1775 => x"00000000",
  1776 => x"00000000",
  1777 => x"00000000",
  1778 => x"00000000",
  1779 => x"00000000",
  1780 => x"00000000",
  1781 => x"00000000",
  1782 => x"00000000",
  1783 => x"00000000",
  1784 => x"00000000",
  1785 => x"00000000",
  1786 => x"00000000",
  1787 => x"00000000",
  1788 => x"00000000",
  1789 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

