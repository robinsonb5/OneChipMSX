-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b0bb5",
     9 => x"ac080b0b",
    10 => x"0bb5b008",
    11 => x"0b0b0bb5",
    12 => x"b4080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"b5b40c0b",
    16 => x"0b0bb5b0",
    17 => x"0c0b0b0b",
    18 => x"b5ac0c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0babf0",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"b5ac70bb",
    57 => x"dc278b38",
    58 => x"80717084",
    59 => x"05530c81",
    60 => x"e2048c51",
    61 => x"8af10402",
    62 => x"fc050df8",
    63 => x"80518f0b",
    64 => x"b5bc0c9f",
    65 => x"0bb5c00c",
    66 => x"a0717081",
    67 => x"055334b5",
    68 => x"c008ff05",
    69 => x"b5c00cb5",
    70 => x"c0088025",
    71 => x"eb38b5bc",
    72 => x"08ff05b5",
    73 => x"bc0cb5bc",
    74 => x"088025d7",
    75 => x"38028405",
    76 => x"0d0402f0",
    77 => x"050df880",
    78 => x"53f8a054",
    79 => x"83bf5273",
    80 => x"70810555",
    81 => x"33517073",
    82 => x"70810555",
    83 => x"34ff1252",
    84 => x"718025eb",
    85 => x"38fbc053",
    86 => x"9f52a073",
    87 => x"70810555",
    88 => x"34ff1252",
    89 => x"718025f2",
    90 => x"38029005",
    91 => x"0d0402f4",
    92 => x"050d7453",
    93 => x"8e0bb5bc",
    94 => x"08258f38",
    95 => x"82b22db5",
    96 => x"bc08ff05",
    97 => x"b5bc0c82",
    98 => x"f404b5bc",
    99 => x"08b5c008",
   100 => x"5351728a",
   101 => x"2e098106",
   102 => x"b7387151",
   103 => x"719f24a0",
   104 => x"38b5bc08",
   105 => x"a02911f8",
   106 => x"80115151",
   107 => x"a07134b5",
   108 => x"c0088105",
   109 => x"b5c00cb5",
   110 => x"c008519f",
   111 => x"7125e238",
   112 => x"800bb5c0",
   113 => x"0cb5bc08",
   114 => x"8105b5bc",
   115 => x"0c83e404",
   116 => x"70a02912",
   117 => x"f8801151",
   118 => x"51727134",
   119 => x"b5c00881",
   120 => x"05b5c00c",
   121 => x"b5c008a0",
   122 => x"2e098106",
   123 => x"8e38800b",
   124 => x"b5c00cb5",
   125 => x"bc088105",
   126 => x"b5bc0c02",
   127 => x"8c050d04",
   128 => x"02e8050d",
   129 => x"77795656",
   130 => x"880bfc16",
   131 => x"77712c8f",
   132 => x"06545254",
   133 => x"80537272",
   134 => x"25953871",
   135 => x"53fbe014",
   136 => x"51877134",
   137 => x"8114ff14",
   138 => x"545472f1",
   139 => x"387153f9",
   140 => x"1576712c",
   141 => x"87065351",
   142 => x"71802e8b",
   143 => x"38fbe014",
   144 => x"51717134",
   145 => x"81145472",
   146 => x"8e249538",
   147 => x"8f733153",
   148 => x"fbe01451",
   149 => x"a0713481",
   150 => x"14ff1454",
   151 => x"5472f138",
   152 => x"0298050d",
   153 => x"0402ec05",
   154 => x"0d800bb5",
   155 => x"c40cf68c",
   156 => x"08f69008",
   157 => x"71882c56",
   158 => x"5481ff06",
   159 => x"52737225",
   160 => x"88387154",
   161 => x"820bb5c4",
   162 => x"0c72882c",
   163 => x"7381ff06",
   164 => x"54557473",
   165 => x"258b3872",
   166 => x"b5c40884",
   167 => x"07b5c40c",
   168 => x"5573842b",
   169 => x"86a07125",
   170 => x"83713170",
   171 => x"0b0b0bb3",
   172 => x"840c8171",
   173 => x"2bff05f6",
   174 => x"880cfecc",
   175 => x"13ff122c",
   176 => x"788829ff",
   177 => x"94057081",
   178 => x"2cb5c408",
   179 => x"52585255",
   180 => x"51525476",
   181 => x"802e8538",
   182 => x"70810751",
   183 => x"70f6940c",
   184 => x"71098105",
   185 => x"f6800c72",
   186 => x"098105f6",
   187 => x"840c0294",
   188 => x"050d0402",
   189 => x"f4050d74",
   190 => x"53727081",
   191 => x"055480f5",
   192 => x"2d527180",
   193 => x"2e893871",
   194 => x"5182ee2d",
   195 => x"85f90402",
   196 => x"8c050d04",
   197 => x"02f8050d",
   198 => x"a5c72d80",
   199 => x"da51a6fe",
   200 => x"2db5ac08",
   201 => x"812a7081",
   202 => x"06515271",
   203 => x"802ee938",
   204 => x"0288050d",
   205 => x"0402f405",
   206 => x"0dbbcc08",
   207 => x"89c406b4",
   208 => x"a00b80f5",
   209 => x"2d525270",
   210 => x"802e8638",
   211 => x"71848007",
   212 => x"52b3d80b",
   213 => x"80f52d72",
   214 => x"07b3f00b",
   215 => x"80f52d70",
   216 => x"812a7081",
   217 => x"06515354",
   218 => x"5270802e",
   219 => x"86387182",
   220 => x"80075272",
   221 => x"81065170",
   222 => x"802e8538",
   223 => x"71880752",
   224 => x"b3fc0b80",
   225 => x"f52d7084",
   226 => x"2b730781",
   227 => x"8432b5ac",
   228 => x"0c51028c",
   229 => x"050d0402",
   230 => x"f4050d74",
   231 => x"70818432",
   232 => x"bbcc0c70",
   233 => x"83065253",
   234 => x"70b3d00b",
   235 => x"880581b7",
   236 => x"2d72892a",
   237 => x"70810651",
   238 => x"5170b4a0",
   239 => x"0b81b72d",
   240 => x"72832a81",
   241 => x"0673882a",
   242 => x"70810651",
   243 => x"52527080",
   244 => x"2e853871",
   245 => x"82075271",
   246 => x"b3f00b81",
   247 => x"b72d7284",
   248 => x"2c708306",
   249 => x"515170b3",
   250 => x"fc0b81b7",
   251 => x"2d70b5ac",
   252 => x"0c028c05",
   253 => x"0d0402d4",
   254 => x"050daec8",
   255 => x"5185f32d",
   256 => x"9c852db5",
   257 => x"ac08802e",
   258 => x"82ab3886",
   259 => x"b52db5ac",
   260 => x"08538ee0",
   261 => x"2db5ac08",
   262 => x"54b5ac08",
   263 => x"802e8297",
   264 => x"389ec82d",
   265 => x"b5ac0880",
   266 => x"2e8738ae",
   267 => x"e05188be",
   268 => x"0497e72d",
   269 => x"b5ac0880",
   270 => x"2e9c38af",
   271 => x"a05185f3",
   272 => x"2d86942d",
   273 => x"72840753",
   274 => x"810bfec4",
   275 => x"0c72fec0",
   276 => x"0c725187",
   277 => x"972d840b",
   278 => x"fec40caf",
   279 => x"e85185f3",
   280 => x"2db08052",
   281 => x"b5cc5194",
   282 => x"fc2db5ac",
   283 => x"089838b0",
   284 => x"8c5185f3",
   285 => x"2db0a452",
   286 => x"b5cc5194",
   287 => x"fc2db5ac",
   288 => x"08802e81",
   289 => x"b038b0b0",
   290 => x"5185f32d",
   291 => x"b5d00857",
   292 => x"8077595a",
   293 => x"767a2e8b",
   294 => x"38811a78",
   295 => x"812a595a",
   296 => x"77f738f7",
   297 => x"1a5a8077",
   298 => x"25818038",
   299 => x"79527751",
   300 => x"84802db5",
   301 => x"d852b5cc",
   302 => x"5197c12d",
   303 => x"b5ac0853",
   304 => x"b5ac0880",
   305 => x"2e80c938",
   306 => x"b5d85b80",
   307 => x"5989fd04",
   308 => x"7a708405",
   309 => x"5c087081",
   310 => x"ff067188",
   311 => x"2c7081ff",
   312 => x"0673902c",
   313 => x"7081ff06",
   314 => x"75982afe",
   315 => x"c80cfec8",
   316 => x"0c58fec8",
   317 => x"0c57fec8",
   318 => x"0c841a5a",
   319 => x"53765384",
   320 => x"80772584",
   321 => x"38848053",
   322 => x"727924c4",
   323 => x"388a9b04",
   324 => x"b0cc5185",
   325 => x"f32d7254",
   326 => x"8ab704b5",
   327 => x"cc519794",
   328 => x"2dfc8017",
   329 => x"81195957",
   330 => x"89a60482",
   331 => x"0bfec40c",
   332 => x"81548ab7",
   333 => x"04805473",
   334 => x"b5ac0c02",
   335 => x"ac050d04",
   336 => x"02f8050d",
   337 => x"a7ce2d81",
   338 => x"f72d8151",
   339 => x"84e52dfe",
   340 => x"c4528172",
   341 => x"0ca58f2d",
   342 => x"a58f2d84",
   343 => x"720c87f6",
   344 => x"2db38851",
   345 => x"a8e72d80",
   346 => x"5184e52d",
   347 => x"0288050d",
   348 => x"0402cc05",
   349 => x"0d8cb851",
   350 => x"87972d81",
   351 => x"0bfec40c",
   352 => x"8cb80bfe",
   353 => x"c00c840b",
   354 => x"fec40c83",
   355 => x"0bfecc0c",
   356 => x"a5aa2da7",
   357 => x"c22da58f",
   358 => x"2da58f2d",
   359 => x"81f72d81",
   360 => x"5184e52d",
   361 => x"a58f2da5",
   362 => x"8f2d8151",
   363 => x"84e52dba",
   364 => x"f451a2d7",
   365 => x"2db5ac08",
   366 => x"ff24f438",
   367 => x"81f452bb",
   368 => x"9c51a39b",
   369 => x"2d87f62d",
   370 => x"b5ac0880",
   371 => x"2e82be38",
   372 => x"8070715b",
   373 => x"585680e4",
   374 => x"76525884",
   375 => x"e52db388",
   376 => x"51a8e72d",
   377 => x"02b40579",
   378 => x"842905f0",
   379 => x"11baf453",
   380 => x"5153a2d7",
   381 => x"2db5ac08",
   382 => x"730cb5ac",
   383 => x"08ff2e09",
   384 => x"81068d38",
   385 => x"ff185877",
   386 => x"80db3877",
   387 => x"598ce504",
   388 => x"81195980",
   389 => x"e4587883",
   390 => x"2e098106",
   391 => x"80c73880",
   392 => x"7a097083",
   393 => x"06fecc0c",
   394 => x"547a7085",
   395 => x"2a708106",
   396 => x"7f585155",
   397 => x"56597279",
   398 => x"2e8a3873",
   399 => x"fe803216",
   400 => x"568cc704",
   401 => x"73165674",
   402 => x"842a7081",
   403 => x"067c5651",
   404 => x"5372802e",
   405 => x"8c387381",
   406 => x"ff321781",
   407 => x"05578ce5",
   408 => x"04767431",
   409 => x"57767607",
   410 => x"5372802e",
   411 => x"80d038fe",
   412 => x"d0087081",
   413 => x"06515372",
   414 => x"802e80c2",
   415 => x"38767655",
   416 => x"5380ff77",
   417 => x"25843880",
   418 => x"ff5380ff",
   419 => x"74258438",
   420 => x"80ff5472",
   421 => x"ff802584",
   422 => x"38ff8053",
   423 => x"73ff8025",
   424 => x"8438ff80",
   425 => x"54767331",
   426 => x"76753174",
   427 => x"882b83fe",
   428 => x"80067681",
   429 => x"ff067107",
   430 => x"fed00c55",
   431 => x"5757a5c7",
   432 => x"2da8f72d",
   433 => x"b5ac0854",
   434 => x"86b52db5",
   435 => x"ac08fec0",
   436 => x"0c86b52d",
   437 => x"b5ac08b5",
   438 => x"c8082e9c",
   439 => x"38b5ac08",
   440 => x"b5c80c84",
   441 => x"53735184",
   442 => x"e52da58f",
   443 => x"2da58f2d",
   444 => x"ff135372",
   445 => x"8025ee38",
   446 => x"73802e89",
   447 => x"388a0bfe",
   448 => x"c40c8be4",
   449 => x"04820bfe",
   450 => x"c40c8be4",
   451 => x"04b0e051",
   452 => x"85f32d82",
   453 => x"0bfec40c",
   454 => x"800bb5ac",
   455 => x"0c02b405",
   456 => x"0d0402e8",
   457 => x"050d7779",
   458 => x"7b585555",
   459 => x"80537276",
   460 => x"25a33874",
   461 => x"70810556",
   462 => x"80f52d74",
   463 => x"70810556",
   464 => x"80f52d52",
   465 => x"5271712e",
   466 => x"86388151",
   467 => x"8ed70481",
   468 => x"13538eae",
   469 => x"04805170",
   470 => x"b5ac0c02",
   471 => x"98050d04",
   472 => x"02d8050d",
   473 => x"800bb9e0",
   474 => x"0cb5d852",
   475 => x"80519da5",
   476 => x"2db5ac08",
   477 => x"54b5ac08",
   478 => x"8c38b0f8",
   479 => x"5185f32d",
   480 => x"73559485",
   481 => x"04805681",
   482 => x"0bba840c",
   483 => x"8853b18c",
   484 => x"52b68e51",
   485 => x"8ea22db5",
   486 => x"ac08762e",
   487 => x"09810687",
   488 => x"38b5ac08",
   489 => x"ba840c88",
   490 => x"53b19852",
   491 => x"b6aa518e",
   492 => x"a22db5ac",
   493 => x"088738b5",
   494 => x"ac08ba84",
   495 => x"0cba8408",
   496 => x"52b1a451",
   497 => x"a0c22dba",
   498 => x"8408802e",
   499 => x"80f638b9",
   500 => x"9e0b80f5",
   501 => x"2db99f0b",
   502 => x"80f52d71",
   503 => x"982b7190",
   504 => x"2b07b9a0",
   505 => x"0b80f52d",
   506 => x"70882b72",
   507 => x"07b9a10b",
   508 => x"80f52d71",
   509 => x"07b9d60b",
   510 => x"80f52db9",
   511 => x"d70b80f5",
   512 => x"2d71882b",
   513 => x"07535f54",
   514 => x"525a5657",
   515 => x"557381ab",
   516 => x"aa2e0981",
   517 => x"068d3875",
   518 => x"519f972d",
   519 => x"b5ac0856",
   520 => x"90b00473",
   521 => x"82d4d52e",
   522 => x"8738b1bc",
   523 => x"5190f104",
   524 => x"b5d85275",
   525 => x"519da52d",
   526 => x"b5ac0855",
   527 => x"b5ac0880",
   528 => x"2e83c238",
   529 => x"8853b198",
   530 => x"52b6aa51",
   531 => x"8ea22db5",
   532 => x"ac088938",
   533 => x"810bb9e0",
   534 => x"0c90f704",
   535 => x"8853b18c",
   536 => x"52b68e51",
   537 => x"8ea22db5",
   538 => x"ac08802e",
   539 => x"8a38b1dc",
   540 => x"5185f32d",
   541 => x"91d104b9",
   542 => x"d60b80f5",
   543 => x"2d547380",
   544 => x"d52e0981",
   545 => x"0680ca38",
   546 => x"b9d70b80",
   547 => x"f52d5473",
   548 => x"81aa2e09",
   549 => x"8106ba38",
   550 => x"800bb5d8",
   551 => x"0b80f52d",
   552 => x"56547481",
   553 => x"e92e8338",
   554 => x"81547481",
   555 => x"eb2e8c38",
   556 => x"80557375",
   557 => x"2e098106",
   558 => x"82cb38b5",
   559 => x"e30b80f5",
   560 => x"2d55748d",
   561 => x"38b5e40b",
   562 => x"80f52d54",
   563 => x"73822e86",
   564 => x"38805594",
   565 => x"8504b5e5",
   566 => x"0b80f52d",
   567 => x"70b9d80c",
   568 => x"ff05b9dc",
   569 => x"0cb5e60b",
   570 => x"80f52db5",
   571 => x"e70b80f5",
   572 => x"2d587605",
   573 => x"77828029",
   574 => x"0570b9e4",
   575 => x"0cb5e80b",
   576 => x"80f52d70",
   577 => x"b9f80cb9",
   578 => x"e0085957",
   579 => x"5876802e",
   580 => x"81a33888",
   581 => x"53b19852",
   582 => x"b6aa518e",
   583 => x"a22db5ac",
   584 => x"0881e238",
   585 => x"b9d80870",
   586 => x"842bb9fc",
   587 => x"0c70b9f4",
   588 => x"0cb5fd0b",
   589 => x"80f52db5",
   590 => x"fc0b80f5",
   591 => x"2d718280",
   592 => x"2905b5fe",
   593 => x"0b80f52d",
   594 => x"70848080",
   595 => x"2912b5ff",
   596 => x"0b80f52d",
   597 => x"7081800a",
   598 => x"291270ba",
   599 => x"800cb9f8",
   600 => x"087129b9",
   601 => x"e4080570",
   602 => x"b9e80cb6",
   603 => x"850b80f5",
   604 => x"2db6840b",
   605 => x"80f52d71",
   606 => x"82802905",
   607 => x"b6860b80",
   608 => x"f52d7084",
   609 => x"80802912",
   610 => x"b6870b80",
   611 => x"f52d7098",
   612 => x"2b81f00a",
   613 => x"06720570",
   614 => x"b9ec0cfe",
   615 => x"117e2977",
   616 => x"05b9f00c",
   617 => x"52595243",
   618 => x"545e5152",
   619 => x"59525d57",
   620 => x"59579483",
   621 => x"04b5ea0b",
   622 => x"80f52db5",
   623 => x"e90b80f5",
   624 => x"2d718280",
   625 => x"290570b9",
   626 => x"fc0c70a0",
   627 => x"2983ff05",
   628 => x"70892a70",
   629 => x"b9f40cb5",
   630 => x"ef0b80f5",
   631 => x"2db5ee0b",
   632 => x"80f52d71",
   633 => x"82802905",
   634 => x"70ba800c",
   635 => x"7b71291e",
   636 => x"70b9f00c",
   637 => x"7db9ec0c",
   638 => x"7305b9e8",
   639 => x"0c555e51",
   640 => x"51555581",
   641 => x"5574b5ac",
   642 => x"0c02a805",
   643 => x"0d0402ec",
   644 => x"050d7670",
   645 => x"872c7180",
   646 => x"ff065556",
   647 => x"54b9e008",
   648 => x"8a387388",
   649 => x"2c7481ff",
   650 => x"065455b5",
   651 => x"d852b9e4",
   652 => x"0815519d",
   653 => x"a52db5ac",
   654 => x"0854b5ac",
   655 => x"08802eb3",
   656 => x"38b9e008",
   657 => x"802e9838",
   658 => x"728429b5",
   659 => x"d8057008",
   660 => x"52539f97",
   661 => x"2db5ac08",
   662 => x"f00a0653",
   663 => x"94f10472",
   664 => x"10b5d805",
   665 => x"7080e02d",
   666 => x"52539fc7",
   667 => x"2db5ac08",
   668 => x"53725473",
   669 => x"b5ac0c02",
   670 => x"94050d04",
   671 => x"02c8050d",
   672 => x"7f615f5b",
   673 => x"800bb9ec",
   674 => x"08b9f008",
   675 => x"595d56b9",
   676 => x"e008762e",
   677 => x"8a38b9d8",
   678 => x"08842b58",
   679 => x"95a504b9",
   680 => x"f408842b",
   681 => x"58805978",
   682 => x"782781a9",
   683 => x"38788f06",
   684 => x"a0175754",
   685 => x"738f38b5",
   686 => x"d8527651",
   687 => x"8117579d",
   688 => x"a52db5d8",
   689 => x"56807680",
   690 => x"f52d5654",
   691 => x"74742e83",
   692 => x"38815474",
   693 => x"81e52e80",
   694 => x"f6388170",
   695 => x"7506555d",
   696 => x"73802e80",
   697 => x"ea388b16",
   698 => x"80f52d98",
   699 => x"065a7980",
   700 => x"de388b53",
   701 => x"7d527551",
   702 => x"8ea22db5",
   703 => x"ac0880cf",
   704 => x"389c1608",
   705 => x"519f972d",
   706 => x"b5ac0884",
   707 => x"1c0c9a16",
   708 => x"80e02d51",
   709 => x"9fc72db5",
   710 => x"ac08b5ac",
   711 => x"08881d0c",
   712 => x"b5ac0855",
   713 => x"55b9e008",
   714 => x"802e9838",
   715 => x"941680e0",
   716 => x"2d519fc7",
   717 => x"2db5ac08",
   718 => x"902b83ff",
   719 => x"f00a0670",
   720 => x"16515473",
   721 => x"881c0c79",
   722 => x"7b0c7c54",
   723 => x"978b0481",
   724 => x"195995a7",
   725 => x"04b9e008",
   726 => x"802eae38",
   727 => x"7b51948e",
   728 => x"2db5ac08",
   729 => x"b5ac0880",
   730 => x"fffffff8",
   731 => x"06555c73",
   732 => x"80ffffff",
   733 => x"f82e9238",
   734 => x"b5ac08fe",
   735 => x"05b9d808",
   736 => x"29b9e808",
   737 => x"055795a5",
   738 => x"04805473",
   739 => x"b5ac0c02",
   740 => x"b8050d04",
   741 => x"02f4050d",
   742 => x"74700881",
   743 => x"05710c70",
   744 => x"08b9dc08",
   745 => x"06535371",
   746 => x"8e388813",
   747 => x"0851948e",
   748 => x"2db5ac08",
   749 => x"88140c81",
   750 => x"0bb5ac0c",
   751 => x"028c050d",
   752 => x"0402f005",
   753 => x"0d758811",
   754 => x"08fe05b9",
   755 => x"d80829b9",
   756 => x"e8081172",
   757 => x"08b9dc08",
   758 => x"06057955",
   759 => x"5354549d",
   760 => x"a52d0290",
   761 => x"050d04b9",
   762 => x"e008b5ac",
   763 => x"0c0402f4",
   764 => x"050dd452",
   765 => x"81ff720c",
   766 => x"71085381",
   767 => x"ff720c72",
   768 => x"882b83fe",
   769 => x"80067208",
   770 => x"7081ff06",
   771 => x"51525381",
   772 => x"ff720c72",
   773 => x"7107882b",
   774 => x"72087081",
   775 => x"ff065152",
   776 => x"5381ff72",
   777 => x"0c727107",
   778 => x"882b7208",
   779 => x"7081ff06",
   780 => x"7207b5ac",
   781 => x"0c525302",
   782 => x"8c050d04",
   783 => x"02f4050d",
   784 => x"74767181",
   785 => x"ff06d40c",
   786 => x"5353ba88",
   787 => x"08853871",
   788 => x"892b5271",
   789 => x"982ad40c",
   790 => x"71902a70",
   791 => x"81ff06d4",
   792 => x"0c517188",
   793 => x"2a7081ff",
   794 => x"06d40c51",
   795 => x"7181ff06",
   796 => x"d40c7290",
   797 => x"2a7081ff",
   798 => x"06d40c51",
   799 => x"d4087081",
   800 => x"ff065151",
   801 => x"82b8bf52",
   802 => x"7081ff2e",
   803 => x"09810694",
   804 => x"3881ff0b",
   805 => x"d40cd408",
   806 => x"7081ff06",
   807 => x"ff145451",
   808 => x"5171e538",
   809 => x"70b5ac0c",
   810 => x"028c050d",
   811 => x"0402fc05",
   812 => x"0d81c751",
   813 => x"81ff0bd4",
   814 => x"0cff1151",
   815 => x"708025f4",
   816 => x"38028405",
   817 => x"0d0402f0",
   818 => x"050d99ad",
   819 => x"2d8fcf53",
   820 => x"805287fc",
   821 => x"80f75198",
   822 => x"bc2db5ac",
   823 => x"0854b5ac",
   824 => x"08812e09",
   825 => x"8106a338",
   826 => x"81ff0bd4",
   827 => x"0c820a52",
   828 => x"849c80e9",
   829 => x"5198bc2d",
   830 => x"b5ac088b",
   831 => x"3881ff0b",
   832 => x"d40c7353",
   833 => x"9a900499",
   834 => x"ad2dff13",
   835 => x"5372c138",
   836 => x"72b5ac0c",
   837 => x"0290050d",
   838 => x"0402f405",
   839 => x"0d81ff0b",
   840 => x"d40c9353",
   841 => x"805287fc",
   842 => x"80c15198",
   843 => x"bc2db5ac",
   844 => x"088b3881",
   845 => x"ff0bd40c",
   846 => x"81539ac6",
   847 => x"0499ad2d",
   848 => x"ff135372",
   849 => x"df3872b5",
   850 => x"ac0c028c",
   851 => x"050d0402",
   852 => x"f0050d99",
   853 => x"ad2d83aa",
   854 => x"52849c80",
   855 => x"c85198bc",
   856 => x"2db5ac08",
   857 => x"812e0981",
   858 => x"06923897",
   859 => x"ee2db5ac",
   860 => x"0883ffff",
   861 => x"06537283",
   862 => x"aa2e9738",
   863 => x"9a992d9b",
   864 => x"8d048154",
   865 => x"9bfc04b1",
   866 => x"fc5185f3",
   867 => x"2d80549b",
   868 => x"fc0481ff",
   869 => x"0bd40cb1",
   870 => x"5399c62d",
   871 => x"b5ac0880",
   872 => x"2e80ca38",
   873 => x"805287fc",
   874 => x"80fa5198",
   875 => x"bc2db5ac",
   876 => x"08b13881",
   877 => x"ff0bd40c",
   878 => x"d4085381",
   879 => x"ff0bd40c",
   880 => x"81ff0bd4",
   881 => x"0c81ff0b",
   882 => x"d40c81ff",
   883 => x"0bd40c72",
   884 => x"862a7081",
   885 => x"06b5ac08",
   886 => x"56515372",
   887 => x"802e9d38",
   888 => x"9b8204b5",
   889 => x"ac0852b2",
   890 => x"9851a0c2",
   891 => x"2d72822e",
   892 => x"ff9538ff",
   893 => x"135372ff",
   894 => x"a0387254",
   895 => x"73b5ac0c",
   896 => x"0290050d",
   897 => x"0402f405",
   898 => x"0d810bba",
   899 => x"880cd008",
   900 => x"708f2a70",
   901 => x"81065151",
   902 => x"5372f338",
   903 => x"72d00c99",
   904 => x"ad2db2a4",
   905 => x"5185f32d",
   906 => x"d008708f",
   907 => x"2a708106",
   908 => x"51515372",
   909 => x"f338810b",
   910 => x"d00c80e3",
   911 => x"53805284",
   912 => x"d480c051",
   913 => x"98bc2db5",
   914 => x"ac08812e",
   915 => x"9a387282",
   916 => x"2e098106",
   917 => x"8c38b2c0",
   918 => x"5185f32d",
   919 => x"80539d9c",
   920 => x"04ff1353",
   921 => x"72d7389a",
   922 => x"cf2db5ac",
   923 => x"08ba880c",
   924 => x"b5ac088b",
   925 => x"38815287",
   926 => x"fc80d051",
   927 => x"98bc2d81",
   928 => x"ff0bd40c",
   929 => x"d008708f",
   930 => x"2a708106",
   931 => x"51515372",
   932 => x"f33872d0",
   933 => x"0c81ff0b",
   934 => x"d40c8153",
   935 => x"72b5ac0c",
   936 => x"028c050d",
   937 => x"0402e005",
   938 => x"0d797b57",
   939 => x"57805881",
   940 => x"ff0bd40c",
   941 => x"d008708f",
   942 => x"2a708106",
   943 => x"51515473",
   944 => x"f3388281",
   945 => x"0bd00c81",
   946 => x"ff0bd40c",
   947 => x"765287fc",
   948 => x"80d15198",
   949 => x"bc2d80db",
   950 => x"c6df55b5",
   951 => x"ac08802e",
   952 => x"9038b5ac",
   953 => x"08537652",
   954 => x"b2d851a0",
   955 => x"c22d9ebf",
   956 => x"0481ff0b",
   957 => x"d40cd408",
   958 => x"7081ff06",
   959 => x"51547381",
   960 => x"fe2e0981",
   961 => x"069d3880",
   962 => x"ff5497ee",
   963 => x"2db5ac08",
   964 => x"76708405",
   965 => x"580cff14",
   966 => x"54738025",
   967 => x"ed388158",
   968 => x"9ea904ff",
   969 => x"155574c9",
   970 => x"3881ff0b",
   971 => x"d40cd008",
   972 => x"708f2a70",
   973 => x"81065151",
   974 => x"5473f338",
   975 => x"73d00c77",
   976 => x"b5ac0c02",
   977 => x"a0050d04",
   978 => x"ba8808b5",
   979 => x"ac0c0402",
   980 => x"e8050d80",
   981 => x"78575575",
   982 => x"70840557",
   983 => x"08538054",
   984 => x"72982a73",
   985 => x"882b5452",
   986 => x"71802ea2",
   987 => x"38c00870",
   988 => x"882a7081",
   989 => x"06515151",
   990 => x"70802ef1",
   991 => x"3871c00c",
   992 => x"81158115",
   993 => x"55558374",
   994 => x"25d63871",
   995 => x"ca3874b5",
   996 => x"ac0c0298",
   997 => x"050d0402",
   998 => x"f4050d74",
   999 => x"70882a83",
  1000 => x"fe800670",
  1001 => x"72982a07",
  1002 => x"72882b87",
  1003 => x"fc808006",
  1004 => x"73982b81",
  1005 => x"f00a0671",
  1006 => x"730707b5",
  1007 => x"ac0c5651",
  1008 => x"5351028c",
  1009 => x"050d0402",
  1010 => x"f8050d02",
  1011 => x"8e0580f5",
  1012 => x"2d74882b",
  1013 => x"077083ff",
  1014 => x"ff06b5ac",
  1015 => x"0c510288",
  1016 => x"050d0402",
  1017 => x"ec050d76",
  1018 => x"53805572",
  1019 => x"75258b38",
  1020 => x"ad5182ee",
  1021 => x"2d720981",
  1022 => x"05537280",
  1023 => x"2eb53887",
  1024 => x"54729c2a",
  1025 => x"73842b54",
  1026 => x"5271802e",
  1027 => x"83388155",
  1028 => x"89722587",
  1029 => x"38b71252",
  1030 => x"a09e04b0",
  1031 => x"12527480",
  1032 => x"2e863871",
  1033 => x"5182ee2d",
  1034 => x"ff145473",
  1035 => x"8025d238",
  1036 => x"a0b804b0",
  1037 => x"5182ee2d",
  1038 => x"800bb5ac",
  1039 => x"0c029405",
  1040 => x"0d0402c0",
  1041 => x"050d0280",
  1042 => x"c4055780",
  1043 => x"70787084",
  1044 => x"055a0872",
  1045 => x"415f5d58",
  1046 => x"7c708405",
  1047 => x"5e085a80",
  1048 => x"5b79982a",
  1049 => x"7a882b5b",
  1050 => x"56758638",
  1051 => x"775fa2ba",
  1052 => x"047d802e",
  1053 => x"81a23880",
  1054 => x"5e7580e4",
  1055 => x"2e8a3875",
  1056 => x"80f82e09",
  1057 => x"81068938",
  1058 => x"76841871",
  1059 => x"085e5854",
  1060 => x"7580e42e",
  1061 => x"9f387580",
  1062 => x"e4268a38",
  1063 => x"7580e32e",
  1064 => x"be38a1ea",
  1065 => x"047580f3",
  1066 => x"2ea33875",
  1067 => x"80f82e89",
  1068 => x"38a1ea04",
  1069 => x"8a53a1bb",
  1070 => x"049053ba",
  1071 => x"8c527b51",
  1072 => x"9fe32db5",
  1073 => x"ac08ba8c",
  1074 => x"5a55a1fa",
  1075 => x"04768418",
  1076 => x"71087054",
  1077 => x"5b58549e",
  1078 => x"cf2d8055",
  1079 => x"a1fa0476",
  1080 => x"84187108",
  1081 => x"585854a2",
  1082 => x"a504a551",
  1083 => x"82ee2d75",
  1084 => x"5182ee2d",
  1085 => x"821858a2",
  1086 => x"ad0474ff",
  1087 => x"16565480",
  1088 => x"7425aa38",
  1089 => x"78708105",
  1090 => x"5a80f52d",
  1091 => x"70525682",
  1092 => x"ee2d8118",
  1093 => x"58a1fa04",
  1094 => x"75a52e09",
  1095 => x"81068638",
  1096 => x"815ea2ad",
  1097 => x"04755182",
  1098 => x"ee2d8118",
  1099 => x"58811b5b",
  1100 => x"837b25fe",
  1101 => x"ac3875fe",
  1102 => x"9f387eb5",
  1103 => x"ac0c0280",
  1104 => x"c0050d04",
  1105 => x"02fc050d",
  1106 => x"72518071",
  1107 => x"0c800b84",
  1108 => x"120c0284",
  1109 => x"050d0402",
  1110 => x"f0050d75",
  1111 => x"70088412",
  1112 => x"08535353",
  1113 => x"ff547171",
  1114 => x"2ea838a7",
  1115 => x"c82d8413",
  1116 => x"08708429",
  1117 => x"14881170",
  1118 => x"087081ff",
  1119 => x"06841808",
  1120 => x"81118706",
  1121 => x"841a0c53",
  1122 => x"51555151",
  1123 => x"51a7c22d",
  1124 => x"715473b5",
  1125 => x"ac0c0290",
  1126 => x"050d0402",
  1127 => x"f4050d74",
  1128 => x"53841308",
  1129 => x"81118706",
  1130 => x"74085451",
  1131 => x"5171712e",
  1132 => x"f038a7c8",
  1133 => x"2d841308",
  1134 => x"70842914",
  1135 => x"88117871",
  1136 => x"0c515151",
  1137 => x"84130881",
  1138 => x"11870684",
  1139 => x"150c51a7",
  1140 => x"c22d028c",
  1141 => x"050d0402",
  1142 => x"f4050da7",
  1143 => x"c82de008",
  1144 => x"e408718b",
  1145 => x"2a708106",
  1146 => x"51535452",
  1147 => x"70802e9d",
  1148 => x"38bacc08",
  1149 => x"708429ba",
  1150 => x"d4057381",
  1151 => x"ff06710c",
  1152 => x"5151bacc",
  1153 => x"08811187",
  1154 => x"06bacc0c",
  1155 => x"51728b2a",
  1156 => x"70810651",
  1157 => x"5170802e",
  1158 => x"b238baf4",
  1159 => x"08708429",
  1160 => x"bafc0574",
  1161 => x"81ff0671",
  1162 => x"0c5151ba",
  1163 => x"f4088111",
  1164 => x"8706baf4",
  1165 => x"0c51baf4",
  1166 => x"08baf808",
  1167 => x"52527171",
  1168 => x"2e098106",
  1169 => x"8638810b",
  1170 => x"bbc40c72",
  1171 => x"8a2a7081",
  1172 => x"06515170",
  1173 => x"802ea838",
  1174 => x"bb9c08bb",
  1175 => x"a0085252",
  1176 => x"71712e9b",
  1177 => x"38bb9c08",
  1178 => x"708429bb",
  1179 => x"a4057008",
  1180 => x"e40c5151",
  1181 => x"bb9c0881",
  1182 => x"118706bb",
  1183 => x"9c0c5180",
  1184 => x"0bbbc80c",
  1185 => x"a7bb2da7",
  1186 => x"c22d028c",
  1187 => x"050d0402",
  1188 => x"fc050da7",
  1189 => x"c82d810b",
  1190 => x"bbc80ca7",
  1191 => x"c22dbbc8",
  1192 => x"085170fa",
  1193 => x"38028405",
  1194 => x"0d0402fc",
  1195 => x"050d800b",
  1196 => x"bbc40cba",
  1197 => x"cc51a2c4",
  1198 => x"2da3d751",
  1199 => x"a7b72da6",
  1200 => x"e12d0284",
  1201 => x"050d0402",
  1202 => x"f4050da6",
  1203 => x"c904b5ac",
  1204 => x"0881f02e",
  1205 => x"09810689",
  1206 => x"38810bb5",
  1207 => x"a00ca6c9",
  1208 => x"04b5ac08",
  1209 => x"81e02e09",
  1210 => x"81068938",
  1211 => x"810bb5a4",
  1212 => x"0ca6c904",
  1213 => x"b5ac0852",
  1214 => x"b5a40880",
  1215 => x"2e8838b5",
  1216 => x"ac088180",
  1217 => x"05527184",
  1218 => x"2c728f06",
  1219 => x"5353b5a0",
  1220 => x"08802e99",
  1221 => x"38728429",
  1222 => x"b4e00572",
  1223 => x"1381712b",
  1224 => x"70097308",
  1225 => x"06730c51",
  1226 => x"5353a6bf",
  1227 => x"04728429",
  1228 => x"b4e00572",
  1229 => x"1383712b",
  1230 => x"72080772",
  1231 => x"0c535380",
  1232 => x"0bb5a40c",
  1233 => x"800bb5a0",
  1234 => x"0cbacc51",
  1235 => x"a2d72db5",
  1236 => x"ac08ff24",
  1237 => x"fef83880",
  1238 => x"0bb5ac0c",
  1239 => x"028c050d",
  1240 => x"0402f805",
  1241 => x"0db4e052",
  1242 => x"8f518072",
  1243 => x"70840554",
  1244 => x"0cff1151",
  1245 => x"708025f2",
  1246 => x"38028805",
  1247 => x"0d0402f0",
  1248 => x"050d7551",
  1249 => x"a7c82d70",
  1250 => x"822cfc06",
  1251 => x"b4e01172",
  1252 => x"109e0671",
  1253 => x"0870722a",
  1254 => x"70830682",
  1255 => x"742b7009",
  1256 => x"7406760c",
  1257 => x"54515657",
  1258 => x"535153a7",
  1259 => x"c22d71b5",
  1260 => x"ac0c0290",
  1261 => x"050d0471",
  1262 => x"980c04ff",
  1263 => x"b008b5ac",
  1264 => x"0c04810b",
  1265 => x"ffb00c04",
  1266 => x"800bffb0",
  1267 => x"0c0402fc",
  1268 => x"050d800b",
  1269 => x"b5a80c80",
  1270 => x"5184e52d",
  1271 => x"0284050d",
  1272 => x"0402f005",
  1273 => x"0dbbd008",
  1274 => x"5481f72d",
  1275 => x"800bbbd4",
  1276 => x"0c730880",
  1277 => x"2e80eb38",
  1278 => x"820bb5c0",
  1279 => x"0cbbd408",
  1280 => x"8f06b5bc",
  1281 => x"0c730852",
  1282 => x"71812ea4",
  1283 => x"3871832e",
  1284 => x"098106b9",
  1285 => x"38881480",
  1286 => x"f52d8415",
  1287 => x"08b2f853",
  1288 => x"545285f3",
  1289 => x"2d718429",
  1290 => x"13700852",
  1291 => x"52a8d104",
  1292 => x"bbcc0888",
  1293 => x"15082c70",
  1294 => x"81065152",
  1295 => x"71802e87",
  1296 => x"38b2fc51",
  1297 => x"a8ca04b3",
  1298 => x"805185f3",
  1299 => x"2d841408",
  1300 => x"5185f32d",
  1301 => x"bbd40881",
  1302 => x"05bbd40c",
  1303 => x"8c1454a7",
  1304 => x"f1040290",
  1305 => x"050d0471",
  1306 => x"bbd00ca7",
  1307 => x"e12dbbd4",
  1308 => x"08ff05bb",
  1309 => x"d80c0402",
  1310 => x"f0050d87",
  1311 => x"51a6fe2d",
  1312 => x"b5ac0881",
  1313 => x"2a708106",
  1314 => x"51527180",
  1315 => x"2ea038a9",
  1316 => x"9504a5c7",
  1317 => x"2d8751a6",
  1318 => x"fe2db5ac",
  1319 => x"08f438b5",
  1320 => x"a8088132",
  1321 => x"70b5a80c",
  1322 => x"70525284",
  1323 => x"e52db5a8",
  1324 => x"08963880",
  1325 => x"da51a6fe",
  1326 => x"2d81f551",
  1327 => x"a6fe2d81",
  1328 => x"f251a6fe",
  1329 => x"2dabe504",
  1330 => x"81f551a6",
  1331 => x"fe2db5ac",
  1332 => x"08812a70",
  1333 => x"81065152",
  1334 => x"71802e8f",
  1335 => x"38bbd808",
  1336 => x"5271802e",
  1337 => x"8638ff12",
  1338 => x"bbd80c81",
  1339 => x"f251a6fe",
  1340 => x"2db5ac08",
  1341 => x"812a7081",
  1342 => x"06515271",
  1343 => x"802e9538",
  1344 => x"bbd408ff",
  1345 => x"05bbd808",
  1346 => x"54527272",
  1347 => x"25863881",
  1348 => x"13bbd80c",
  1349 => x"80da51a6",
  1350 => x"fe2db5ac",
  1351 => x"08812a70",
  1352 => x"81065152",
  1353 => x"71802e80",
  1354 => x"fb38bbd0",
  1355 => x"08bbd808",
  1356 => x"55537380",
  1357 => x"2e8a388c",
  1358 => x"13ff1555",
  1359 => x"53aab204",
  1360 => x"72085271",
  1361 => x"822ea638",
  1362 => x"71822689",
  1363 => x"3871812e",
  1364 => x"a538aba4",
  1365 => x"0471832e",
  1366 => x"ad387184",
  1367 => x"2e098106",
  1368 => x"80c23888",
  1369 => x"130851a8",
  1370 => x"e72daba4",
  1371 => x"04881308",
  1372 => x"52712dab",
  1373 => x"a404810b",
  1374 => x"8814082b",
  1375 => x"bbcc0832",
  1376 => x"bbcc0cab",
  1377 => x"a1048813",
  1378 => x"80f52d81",
  1379 => x"058b1480",
  1380 => x"f52d5354",
  1381 => x"71742483",
  1382 => x"38805473",
  1383 => x"881481b7",
  1384 => x"2da7e12d",
  1385 => x"8054800b",
  1386 => x"b5c00c73",
  1387 => x"8f06b5bc",
  1388 => x"0ca05273",
  1389 => x"bbd8082e",
  1390 => x"09810698",
  1391 => x"38bbd408",
  1392 => x"ff057432",
  1393 => x"70098105",
  1394 => x"7072079f",
  1395 => x"2a917131",
  1396 => x"51515353",
  1397 => x"715182ee",
  1398 => x"2d811454",
  1399 => x"8e7425c6",
  1400 => x"38b5a808",
  1401 => x"5271b5ac",
  1402 => x"0c029005",
  1403 => x"0d040000",
  1404 => x"00ffffff",
  1405 => x"ff00ffff",
  1406 => x"ffff00ff",
  1407 => x"ffffff00",
  1408 => x"52657365",
  1409 => x"74000000",
  1410 => x"4f707469",
  1411 => x"6f6e7320",
  1412 => x"10000000",
  1413 => x"54757262",
  1414 => x"6f202831",
  1415 => x"302e3734",
  1416 => x"4d487a29",
  1417 => x"00000000",
  1418 => x"4d6f7573",
  1419 => x"6520656d",
  1420 => x"756c6174",
  1421 => x"696f6e00",
  1422 => x"45786974",
  1423 => x"00000000",
  1424 => x"53442043",
  1425 => x"61726400",
  1426 => x"4a617061",
  1427 => x"6e657365",
  1428 => x"206b6579",
  1429 => x"626f6172",
  1430 => x"64206c61",
  1431 => x"796f7574",
  1432 => x"00000000",
  1433 => x"4261636b",
  1434 => x"00000000",
  1435 => x"32303438",
  1436 => x"4c422052",
  1437 => x"414d0000",
  1438 => x"34303936",
  1439 => x"4b422052",
  1440 => x"414d0000",
  1441 => x"536c323a",
  1442 => x"204e6f6e",
  1443 => x"65000000",
  1444 => x"536c323a",
  1445 => x"20455345",
  1446 => x"2d534343",
  1447 => x"20314d42",
  1448 => x"2f534343",
  1449 => x"2d490000",
  1450 => x"536c323a",
  1451 => x"20455345",
  1452 => x"2d52414d",
  1453 => x"20314d42",
  1454 => x"2f415343",
  1455 => x"49493800",
  1456 => x"536c323a",
  1457 => x"20455345",
  1458 => x"2d52414d",
  1459 => x"20314d42",
  1460 => x"2f415343",
  1461 => x"49493136",
  1462 => x"00000000",
  1463 => x"536c313a",
  1464 => x"204e6f6e",
  1465 => x"65000000",
  1466 => x"536c313a",
  1467 => x"20455345",
  1468 => x"2d534343",
  1469 => x"20314d42",
  1470 => x"2f534343",
  1471 => x"2d490000",
  1472 => x"536c313a",
  1473 => x"204d6567",
  1474 => x"6152414d",
  1475 => x"00000000",
  1476 => x"56474120",
  1477 => x"2d203331",
  1478 => x"4b487a2c",
  1479 => x"20363048",
  1480 => x"7a000000",
  1481 => x"56474120",
  1482 => x"2d203331",
  1483 => x"4b487a2c",
  1484 => x"20353048",
  1485 => x"7a000000",
  1486 => x"5456202d",
  1487 => x"20343830",
  1488 => x"692c2036",
  1489 => x"30487a00",
  1490 => x"496e6974",
  1491 => x"69616c69",
  1492 => x"7a696e67",
  1493 => x"20534420",
  1494 => x"63617264",
  1495 => x"0a000000",
  1496 => x"53444843",
  1497 => x"20636172",
  1498 => x"64206465",
  1499 => x"74656374",
  1500 => x"65642062",
  1501 => x"7574206e",
  1502 => x"6f740a73",
  1503 => x"7570706f",
  1504 => x"72746564",
  1505 => x"3b206469",
  1506 => x"7361626c",
  1507 => x"696e6720",
  1508 => x"53442063",
  1509 => x"6172640a",
  1510 => x"10204f4b",
  1511 => x"0a000000",
  1512 => x"46617433",
  1513 => x"32206669",
  1514 => x"6c657379",
  1515 => x"7374656d",
  1516 => x"20646574",
  1517 => x"65637465",
  1518 => x"64206275",
  1519 => x"740a6e6f",
  1520 => x"74207375",
  1521 => x"70706f72",
  1522 => x"7465643b",
  1523 => x"20646973",
  1524 => x"61626c69",
  1525 => x"6e672053",
  1526 => x"44206361",
  1527 => x"72640a10",
  1528 => x"204f4b0a",
  1529 => x"00000000",
  1530 => x"54727969",
  1531 => x"6e67204d",
  1532 => x"53583342",
  1533 => x"494f532e",
  1534 => x"5359532e",
  1535 => x"2e2e0a00",
  1536 => x"4d535833",
  1537 => x"42494f53",
  1538 => x"53595300",
  1539 => x"54727969",
  1540 => x"6e672042",
  1541 => x"494f535f",
  1542 => x"4d32502e",
  1543 => x"524f4d2e",
  1544 => x"2e2e0a00",
  1545 => x"42494f53",
  1546 => x"5f4d3250",
  1547 => x"524f4d00",
  1548 => x"4f70656e",
  1549 => x"65642042",
  1550 => x"494f532c",
  1551 => x"206c6f61",
  1552 => x"64696e67",
  1553 => x"2e2e2e0a",
  1554 => x"00000000",
  1555 => x"52656164",
  1556 => x"20626c6f",
  1557 => x"636b2066",
  1558 => x"61696c65",
  1559 => x"640a0000",
  1560 => x"4c6f6164",
  1561 => x"696e6720",
  1562 => x"42494f53",
  1563 => x"20666169",
  1564 => x"6c65640a",
  1565 => x"00000000",
  1566 => x"52656164",
  1567 => x"206f6620",
  1568 => x"4d425220",
  1569 => x"6661696c",
  1570 => x"65640a00",
  1571 => x"46415431",
  1572 => x"36202020",
  1573 => x"00000000",
  1574 => x"46415433",
  1575 => x"32202020",
  1576 => x"00000000",
  1577 => x"25642070",
  1578 => x"61727469",
  1579 => x"74696f6e",
  1580 => x"7320666f",
  1581 => x"756e640a",
  1582 => x"00000000",
  1583 => x"4e6f2070",
  1584 => x"61727469",
  1585 => x"74696f6e",
  1586 => x"20736967",
  1587 => x"6e617475",
  1588 => x"72652066",
  1589 => x"6f756e64",
  1590 => x"0a000000",
  1591 => x"556e7375",
  1592 => x"70706f72",
  1593 => x"74656420",
  1594 => x"70617274",
  1595 => x"6974696f",
  1596 => x"6e207479",
  1597 => x"7065210a",
  1598 => x"00000000",
  1599 => x"53444843",
  1600 => x"20496e69",
  1601 => x"7469616c",
  1602 => x"697a6174",
  1603 => x"696f6e20",
  1604 => x"6572726f",
  1605 => x"72210a00",
  1606 => x"434d4435",
  1607 => x"38202564",
  1608 => x"0a202000",
  1609 => x"496e6974",
  1610 => x"69616c69",
  1611 => x"7a696e67",
  1612 => x"20534420",
  1613 => x"63617264",
  1614 => x"2e2e2e0a",
  1615 => x"00000000",
  1616 => x"53442063",
  1617 => x"61726420",
  1618 => x"72657365",
  1619 => x"74206661",
  1620 => x"696c6564",
  1621 => x"210a0000",
  1622 => x"52656164",
  1623 => x"20636f6d",
  1624 => x"6d616e64",
  1625 => x"20666169",
  1626 => x"6c656420",
  1627 => x"61742025",
  1628 => x"64202825",
  1629 => x"64290a00",
  1630 => x"16200000",
  1631 => x"14200000",
  1632 => x"15200000",
  1633 => x"00000002",
  1634 => x"00000002",
  1635 => x"00001600",
  1636 => x"00000540",
  1637 => x"00000004",
  1638 => x"00001608",
  1639 => x"000019d0",
  1640 => x"00000001",
  1641 => x"00001614",
  1642 => x"00000007",
  1643 => x"00000001",
  1644 => x"00001628",
  1645 => x"0000000a",
  1646 => x"00000002",
  1647 => x"00001638",
  1648 => x"000013ce",
  1649 => x"00000000",
  1650 => x"00000000",
  1651 => x"00000000",
  1652 => x"00000003",
  1653 => x"00001a54",
  1654 => x"00000003",
  1655 => x"00000001",
  1656 => x"00001640",
  1657 => x"00000002",
  1658 => x"00000003",
  1659 => x"00001a48",
  1660 => x"00000003",
  1661 => x"00000003",
  1662 => x"00001a38",
  1663 => x"00000004",
  1664 => x"00000001",
  1665 => x"00001648",
  1666 => x"00000006",
  1667 => x"00000003",
  1668 => x"00001a30",
  1669 => x"00000002",
  1670 => x"00000004",
  1671 => x"00001664",
  1672 => x"00001988",
  1673 => x"00000000",
  1674 => x"00000000",
  1675 => x"00000000",
  1676 => x"0000166c",
  1677 => x"00001678",
  1678 => x"00001684",
  1679 => x"00001690",
  1680 => x"000016a8",
  1681 => x"000016c0",
  1682 => x"000016dc",
  1683 => x"000016e8",
  1684 => x"00001700",
  1685 => x"00001710",
  1686 => x"00001724",
  1687 => x"00001738",
  1688 => x"00000000",
  1689 => x"00000000",
  1690 => x"00000000",
  1691 => x"00000000",
  1692 => x"00000000",
  1693 => x"00000000",
  1694 => x"00000000",
  1695 => x"00000000",
  1696 => x"00000000",
  1697 => x"00000000",
  1698 => x"00000000",
  1699 => x"00000000",
  1700 => x"00000000",
  1701 => x"00000000",
  1702 => x"00000000",
  1703 => x"00000000",
  1704 => x"00000000",
  1705 => x"00000000",
  1706 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

