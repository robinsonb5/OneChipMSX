-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b0bb3",
     9 => x"e4080b0b",
    10 => x"0bb3e808",
    11 => x"0b0b0bb3",
    12 => x"ec080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"b3ec0c0b",
    16 => x"0b0bb3e8",
    17 => x"0c0b0b0b",
    18 => x"b3e40c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0ba490",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"b3e470ba",
    57 => x"bc278b38",
    58 => x"80717084",
    59 => x"05530c81",
    60 => x"e2048c51",
    61 => x"81f70402",
    62 => x"d8050d81",
    63 => x"0bfec40c",
    64 => x"b90bfec0",
    65 => x"0c840bfe",
    66 => x"c40ca4a0",
    67 => x"5195d32d",
    68 => x"9efc2da2",
    69 => x"aa2da4c0",
    70 => x"5195d32d",
    71 => x"92ef2db3",
    72 => x"e408802e",
    73 => x"81c538a4",
    74 => x"d85195d3",
    75 => x"2d84c22d",
    76 => x"a4f052b5",
    77 => x"9c518b97",
    78 => x"2db3e408",
    79 => x"81ff0653",
    80 => x"72802e81",
    81 => x"a038a4fc",
    82 => x"5195d32d",
    83 => x"b5a00857",
    84 => x"80597877",
    85 => x"25819438",
    86 => x"b5b452b5",
    87 => x"9c518dee",
    88 => x"2db3e408",
    89 => x"81ff06b5",
    90 => x"b45b5380",
    91 => x"5872782e",
    92 => x"098106b1",
    93 => x"3883b804",
    94 => x"79708405",
    95 => x"5b087081",
    96 => x"ff067188",
    97 => x"2c7081ff",
    98 => x"0673902c",
    99 => x"7081ff06",
   100 => x"75982afe",
   101 => x"c80cfec8",
   102 => x"0c58fec8",
   103 => x"0c57fec8",
   104 => x"0c841959",
   105 => x"53765384",
   106 => x"80772584",
   107 => x"38848053",
   108 => x"727824c4",
   109 => x"3883be04",
   110 => x"a5985195",
   111 => x"d32db59c",
   112 => x"518dc12d",
   113 => x"fc801781",
   114 => x"1a5a57ae",
   115 => x"5195b12d",
   116 => x"78bf0653",
   117 => x"7286388a",
   118 => x"5195b12d",
   119 => x"768024fe",
   120 => x"f73883eb",
   121 => x"04a5ac51",
   122 => x"95d32d82",
   123 => x"0bfec40c",
   124 => x"9f942db3",
   125 => x"e408802e",
   126 => x"f738b3e4",
   127 => x"085195b1",
   128 => x"2d83f004",
   129 => x"02e8050d",
   130 => x"77797b58",
   131 => x"55558053",
   132 => x"727625a3",
   133 => x"38747081",
   134 => x"055680f5",
   135 => x"2d747081",
   136 => x"055680f5",
   137 => x"2d525271",
   138 => x"712e8638",
   139 => x"815184b9",
   140 => x"04811353",
   141 => x"84900480",
   142 => x"5170b3e4",
   143 => x"0c029805",
   144 => x"0d0402d8",
   145 => x"050d800b",
   146 => x"b9cc0ca5",
   147 => x"c45195d3",
   148 => x"2db5b452",
   149 => x"8051948e",
   150 => x"2db3e408",
   151 => x"54b3e408",
   152 => x"8c38a5d4",
   153 => x"5195d32d",
   154 => x"73558a95",
   155 => x"04a5e851",
   156 => x"95d32d80",
   157 => x"56810bb5",
   158 => x"a80c8853",
   159 => x"a68052b5",
   160 => x"ea518484",
   161 => x"2db3e408",
   162 => x"762e0981",
   163 => x"068738b3",
   164 => x"e408b5a8",
   165 => x"0c8853a6",
   166 => x"8c52b686",
   167 => x"5184842d",
   168 => x"b3e40887",
   169 => x"38b3e408",
   170 => x"b5a80cb5",
   171 => x"a80852a6",
   172 => x"985197db",
   173 => x"2db5a808",
   174 => x"802e8187",
   175 => x"38b8fa0b",
   176 => x"80f52db8",
   177 => x"fb0b80f5",
   178 => x"2d71982b",
   179 => x"71902b07",
   180 => x"b8fc0b80",
   181 => x"f52d7088",
   182 => x"2b7207b8",
   183 => x"fd0b80f5",
   184 => x"2d7107b9",
   185 => x"b20b80f5",
   186 => x"2db9b30b",
   187 => x"80f52d71",
   188 => x"882b0753",
   189 => x"5f54525a",
   190 => x"56575573",
   191 => x"81abaa2e",
   192 => x"0981068d",
   193 => x"38755196",
   194 => x"9b2db3e4",
   195 => x"085686a1",
   196 => x"047382d4",
   197 => x"d52e8a38",
   198 => x"a6ac5195",
   199 => x"d32d87d6",
   200 => x"047552a6",
   201 => x"cc5197db",
   202 => x"2db5b452",
   203 => x"7551948e",
   204 => x"2db3e408",
   205 => x"55b3e408",
   206 => x"802e83d9",
   207 => x"38a6e451",
   208 => x"95d32da7",
   209 => x"8c5197db",
   210 => x"2d8853a6",
   211 => x"8c52b686",
   212 => x"5184842d",
   213 => x"b3e40889",
   214 => x"38810bb9",
   215 => x"cc0c86fc",
   216 => x"048853a6",
   217 => x"8052b5ea",
   218 => x"5184842d",
   219 => x"b3e40880",
   220 => x"2e8a38a7",
   221 => x"a45197db",
   222 => x"2d87d604",
   223 => x"b9b20b80",
   224 => x"f52d5473",
   225 => x"80d52e09",
   226 => x"810680ca",
   227 => x"38b9b30b",
   228 => x"80f52d54",
   229 => x"7381aa2e",
   230 => x"098106ba",
   231 => x"38800bb5",
   232 => x"b40b80f5",
   233 => x"2d565474",
   234 => x"81e92e83",
   235 => x"38815474",
   236 => x"81eb2e8c",
   237 => x"38805573",
   238 => x"752e0981",
   239 => x"0682d638",
   240 => x"b5bf0b80",
   241 => x"f52d5978",
   242 => x"8d38b5c0",
   243 => x"0b80f52d",
   244 => x"5473822e",
   245 => x"86388055",
   246 => x"8a9504b5",
   247 => x"c10b80f5",
   248 => x"2d70b9d4",
   249 => x"0cff1170",
   250 => x"b9c80c54",
   251 => x"52a7c451",
   252 => x"97db2db5",
   253 => x"c20b80f5",
   254 => x"2db5c30b",
   255 => x"80f52d56",
   256 => x"76057582",
   257 => x"80290570",
   258 => x"b9bc0cb5",
   259 => x"c40b80f5",
   260 => x"2d70b9b8",
   261 => x"0cb9cc08",
   262 => x"59575876",
   263 => x"802e81a5",
   264 => x"388853a6",
   265 => x"8c52b686",
   266 => x"5184842d",
   267 => x"7855b3e4",
   268 => x"0881e238",
   269 => x"b9d40870",
   270 => x"842bb9b4",
   271 => x"0c70b9d0",
   272 => x"0cb5d90b",
   273 => x"80f52db5",
   274 => x"d80b80f5",
   275 => x"2d718280",
   276 => x"2905b5da",
   277 => x"0b80f52d",
   278 => x"70848080",
   279 => x"2912b5db",
   280 => x"0b80f52d",
   281 => x"7081800a",
   282 => x"291270b5",
   283 => x"ac0cb9b8",
   284 => x"087129b9",
   285 => x"bc080570",
   286 => x"b9dc0cb5",
   287 => x"e10b80f5",
   288 => x"2db5e00b",
   289 => x"80f52d71",
   290 => x"82802905",
   291 => x"b5e20b80",
   292 => x"f52d7084",
   293 => x"80802912",
   294 => x"b5e30b80",
   295 => x"f52d7098",
   296 => x"2b81f00a",
   297 => x"06720570",
   298 => x"b5b00cfe",
   299 => x"117e2977",
   300 => x"05b9c40c",
   301 => x"52575257",
   302 => x"5d575152",
   303 => x"5f525c57",
   304 => x"57578a93",
   305 => x"04b5c60b",
   306 => x"80f52db5",
   307 => x"c50b80f5",
   308 => x"2d718280",
   309 => x"290570b9",
   310 => x"b40c70a0",
   311 => x"2983ff05",
   312 => x"70892a70",
   313 => x"b9d00cb5",
   314 => x"cb0b80f5",
   315 => x"2db5ca0b",
   316 => x"80f52d71",
   317 => x"82802905",
   318 => x"70b5ac0c",
   319 => x"7b71291e",
   320 => x"70b9c40c",
   321 => x"7db5b00c",
   322 => x"7305b9dc",
   323 => x"0c555e51",
   324 => x"51555581",
   325 => x"5574b3e4",
   326 => x"0c02a805",
   327 => x"0d0402ec",
   328 => x"050d7670",
   329 => x"872c7180",
   330 => x"ff065755",
   331 => x"53b9cc08",
   332 => x"8a387288",
   333 => x"2c7381ff",
   334 => x"065654b9",
   335 => x"bc081452",
   336 => x"a7e85197",
   337 => x"db2db5b4",
   338 => x"52b9bc08",
   339 => x"1451948e",
   340 => x"2db3e408",
   341 => x"53b3e408",
   342 => x"802eb338",
   343 => x"b9cc0880",
   344 => x"2e983874",
   345 => x"8429b5b4",
   346 => x"05700852",
   347 => x"53969b2d",
   348 => x"b3e408f0",
   349 => x"0a06558b",
   350 => x"8c047410",
   351 => x"b5b40570",
   352 => x"80e02d52",
   353 => x"5396cb2d",
   354 => x"b3e40855",
   355 => x"745372b3",
   356 => x"e40c0294",
   357 => x"050d0402",
   358 => x"c8050d7f",
   359 => x"615f5c80",
   360 => x"0bb5b008",
   361 => x"b9c40859",
   362 => x"5956b9cc",
   363 => x"08762e8a",
   364 => x"38b9d408",
   365 => x"842b598b",
   366 => x"c004b9d0",
   367 => x"08842b59",
   368 => x"805a7979",
   369 => x"2781b638",
   370 => x"798f06a0",
   371 => x"17575473",
   372 => x"97387652",
   373 => x"a8885197",
   374 => x"db2db5b4",
   375 => x"52765181",
   376 => x"1757948e",
   377 => x"2db5b456",
   378 => x"807680f5",
   379 => x"2d565474",
   380 => x"742e8338",
   381 => x"81547481",
   382 => x"e52e80fb",
   383 => x"38817075",
   384 => x"06555d73",
   385 => x"802e80ef",
   386 => x"388b1680",
   387 => x"f52d9806",
   388 => x"5b7a80e3",
   389 => x"38755195",
   390 => x"d32d8b53",
   391 => x"7d527551",
   392 => x"84842db3",
   393 => x"e40880cf",
   394 => x"389c1608",
   395 => x"51969b2d",
   396 => x"b3e40884",
   397 => x"1d0c9a16",
   398 => x"80e02d51",
   399 => x"96cb2db3",
   400 => x"e408b3e4",
   401 => x"08881e0c",
   402 => x"b3e40855",
   403 => x"55b9cc08",
   404 => x"802e9838",
   405 => x"941680e0",
   406 => x"2d5196cb",
   407 => x"2db3e408",
   408 => x"902b83ff",
   409 => x"f00a0670",
   410 => x"16515473",
   411 => x"881d0c7a",
   412 => x"7c0c7c54",
   413 => x"8db80481",
   414 => x"1a5a8bc2",
   415 => x"04b9cc08",
   416 => x"802eb338",
   417 => x"77518a9e",
   418 => x"2db3e408",
   419 => x"b3e40853",
   420 => x"a8a85258",
   421 => x"97db2d77",
   422 => x"80ffffff",
   423 => x"f8065473",
   424 => x"80ffffff",
   425 => x"f82e8f38",
   426 => x"fe18b9d4",
   427 => x"0829b9dc",
   428 => x"0805578b",
   429 => x"c0048054",
   430 => x"73b3e40c",
   431 => x"02b8050d",
   432 => x"0402f405",
   433 => x"0d747008",
   434 => x"8105710c",
   435 => x"7008b9c8",
   436 => x"08065353",
   437 => x"718e3888",
   438 => x"1308518a",
   439 => x"9e2db3e4",
   440 => x"0888140c",
   441 => x"810bb3e4",
   442 => x"0c028c05",
   443 => x"0d0402f0",
   444 => x"050d7588",
   445 => x"1108fe05",
   446 => x"b9d40829",
   447 => x"b9dc0811",
   448 => x"7208b9c8",
   449 => x"08060579",
   450 => x"55535454",
   451 => x"948e2db3",
   452 => x"e40853b3",
   453 => x"e408802e",
   454 => x"83388153",
   455 => x"72b3e40c",
   456 => x"0290050d",
   457 => x"0402f405",
   458 => x"0dd45281",
   459 => x"ff720c71",
   460 => x"085381ff",
   461 => x"720c7288",
   462 => x"2b83fe80",
   463 => x"06720870",
   464 => x"81ff0651",
   465 => x"525381ff",
   466 => x"720c7271",
   467 => x"07882b72",
   468 => x"087081ff",
   469 => x"06515253",
   470 => x"81ff720c",
   471 => x"72710788",
   472 => x"2b720870",
   473 => x"81ff0672",
   474 => x"07b3e40c",
   475 => x"5253028c",
   476 => x"050d0402",
   477 => x"f4050d74",
   478 => x"767181ff",
   479 => x"06d40c53",
   480 => x"53b9e008",
   481 => x"85387189",
   482 => x"2b527198",
   483 => x"2ad40c71",
   484 => x"902a7081",
   485 => x"ff06d40c",
   486 => x"5171882a",
   487 => x"7081ff06",
   488 => x"d40c5171",
   489 => x"81ff06d4",
   490 => x"0c72902a",
   491 => x"7081ff06",
   492 => x"d40c51d4",
   493 => x"087081ff",
   494 => x"06515182",
   495 => x"b8bf5270",
   496 => x"81ff2e09",
   497 => x"81069438",
   498 => x"81ff0bd4",
   499 => x"0cd40870",
   500 => x"81ff06ff",
   501 => x"14545151",
   502 => x"71e53870",
   503 => x"b3e40c02",
   504 => x"8c050d04",
   505 => x"02fc050d",
   506 => x"81c75181",
   507 => x"ff0bd40c",
   508 => x"ff115170",
   509 => x"8025f438",
   510 => x"0284050d",
   511 => x"0402f005",
   512 => x"0d8fe42d",
   513 => x"819c9f53",
   514 => x"805287fc",
   515 => x"80f7518e",
   516 => x"f32db3e4",
   517 => x"0854b3e4",
   518 => x"08812e09",
   519 => x"8106a338",
   520 => x"81ff0bd4",
   521 => x"0c820a52",
   522 => x"849c80e9",
   523 => x"518ef32d",
   524 => x"b3e4088b",
   525 => x"3881ff0b",
   526 => x"d40c7353",
   527 => x"90c8048f",
   528 => x"e42dff13",
   529 => x"5372c138",
   530 => x"72b3e40c",
   531 => x"0290050d",
   532 => x"0402f405",
   533 => x"0d81ff0b",
   534 => x"d40ca8c0",
   535 => x"5195d32d",
   536 => x"93538052",
   537 => x"87fc80c1",
   538 => x"518ef32d",
   539 => x"b3e4088b",
   540 => x"3881ff0b",
   541 => x"d40c8153",
   542 => x"9184048f",
   543 => x"e42dff13",
   544 => x"5372df38",
   545 => x"72b3e40c",
   546 => x"028c050d",
   547 => x"0402f005",
   548 => x"0d8fe42d",
   549 => x"83aa5284",
   550 => x"9c80c851",
   551 => x"8ef32db3",
   552 => x"e408b3e4",
   553 => x"0853a8cc",
   554 => x"525397db",
   555 => x"2d72812e",
   556 => x"0981069c",
   557 => x"388ea52d",
   558 => x"b3e40883",
   559 => x"ffff0653",
   560 => x"7283aa2e",
   561 => x"a138b3e4",
   562 => x"0852a8e4",
   563 => x"5197db2d",
   564 => x"90d12d91",
   565 => x"e1048154",
   566 => x"92e604a8",
   567 => x"fc5197db",
   568 => x"2d805492",
   569 => x"e60481ff",
   570 => x"0bd40cb1",
   571 => x"538ffd2d",
   572 => x"b3e40880",
   573 => x"2e80e038",
   574 => x"805287fc",
   575 => x"80fa518e",
   576 => x"f32db3e4",
   577 => x"0880c638",
   578 => x"b3e40852",
   579 => x"a9985197",
   580 => x"db2d81ff",
   581 => x"0bd40cd4",
   582 => x"087081ff",
   583 => x"067054a9",
   584 => x"a4535153",
   585 => x"97db2d81",
   586 => x"ff0bd40c",
   587 => x"81ff0bd4",
   588 => x"0c81ff0b",
   589 => x"d40c81ff",
   590 => x"0bd40c72",
   591 => x"862a7081",
   592 => x"06705651",
   593 => x"5372802e",
   594 => x"9d3891d6",
   595 => x"04b3e408",
   596 => x"52a99851",
   597 => x"97db2d72",
   598 => x"822efeff",
   599 => x"38ff1353",
   600 => x"72ff8a38",
   601 => x"725473b3",
   602 => x"e40c0290",
   603 => x"050d0402",
   604 => x"f4050d81",
   605 => x"0bb9e00c",
   606 => x"d008708f",
   607 => x"2a708106",
   608 => x"51515372",
   609 => x"f33872d0",
   610 => x"0c8fe42d",
   611 => x"a9b45195",
   612 => x"d32dd008",
   613 => x"708f2a70",
   614 => x"81065151",
   615 => x"5372f338",
   616 => x"810bd00c",
   617 => x"87538052",
   618 => x"84d480c0",
   619 => x"518ef32d",
   620 => x"b3e40881",
   621 => x"2e943872",
   622 => x"822e0981",
   623 => x"06863880",
   624 => x"5393ff04",
   625 => x"ff135372",
   626 => x"dd38918d",
   627 => x"2db3e408",
   628 => x"b9e00cb3",
   629 => x"e4088b38",
   630 => x"815287fc",
   631 => x"80d0518e",
   632 => x"f32d81ff",
   633 => x"0bd40cd0",
   634 => x"08708f2a",
   635 => x"70810651",
   636 => x"515372f3",
   637 => x"3872d00c",
   638 => x"81ff0bd4",
   639 => x"0c815372",
   640 => x"b3e40c02",
   641 => x"8c050d04",
   642 => x"800bb3e4",
   643 => x"0c0402e0",
   644 => x"050d797b",
   645 => x"57578058",
   646 => x"81ff0bd4",
   647 => x"0cd00870",
   648 => x"8f2a7081",
   649 => x"06515154",
   650 => x"73f33882",
   651 => x"810bd00c",
   652 => x"81ff0bd4",
   653 => x"0c765287",
   654 => x"fc80d151",
   655 => x"8ef32d80",
   656 => x"dbc6df55",
   657 => x"b3e40880",
   658 => x"2e9038b3",
   659 => x"e4085376",
   660 => x"52a9c051",
   661 => x"97db2d95",
   662 => x"a80481ff",
   663 => x"0bd40cd4",
   664 => x"087081ff",
   665 => x"06515473",
   666 => x"81fe2e09",
   667 => x"81069d38",
   668 => x"80ff548e",
   669 => x"a52db3e4",
   670 => x"08767084",
   671 => x"05580cff",
   672 => x"14547380",
   673 => x"25ed3881",
   674 => x"58959204",
   675 => x"ff155574",
   676 => x"c93881ff",
   677 => x"0bd40cd0",
   678 => x"08708f2a",
   679 => x"70810651",
   680 => x"515473f3",
   681 => x"3873d00c",
   682 => x"77b3e40c",
   683 => x"02a0050d",
   684 => x"0402f805",
   685 => x"0d7352c0",
   686 => x"0870882a",
   687 => x"70810651",
   688 => x"51517080",
   689 => x"2ef13871",
   690 => x"c00c71b3",
   691 => x"e40c0288",
   692 => x"050d0402",
   693 => x"e8050d80",
   694 => x"78575575",
   695 => x"70840557",
   696 => x"08538054",
   697 => x"72982a73",
   698 => x"882b5452",
   699 => x"71802ea2",
   700 => x"38c00870",
   701 => x"882a7081",
   702 => x"06515151",
   703 => x"70802ef1",
   704 => x"3871c00c",
   705 => x"81158115",
   706 => x"55558374",
   707 => x"25d63871",
   708 => x"ca3874b3",
   709 => x"e40c0298",
   710 => x"050d0402",
   711 => x"f4050d74",
   712 => x"70882a83",
   713 => x"fe800670",
   714 => x"72982a07",
   715 => x"72882b87",
   716 => x"fc808006",
   717 => x"73982b81",
   718 => x"f00a0671",
   719 => x"730707b3",
   720 => x"e40c5651",
   721 => x"5351028c",
   722 => x"050d0402",
   723 => x"f8050d02",
   724 => x"8e0580f5",
   725 => x"2d74882b",
   726 => x"077083ff",
   727 => x"ff06b3e4",
   728 => x"0c510288",
   729 => x"050d0402",
   730 => x"f8050d73",
   731 => x"70902b71",
   732 => x"902a07b3",
   733 => x"e40c5202",
   734 => x"88050d04",
   735 => x"02ec050d",
   736 => x"76538055",
   737 => x"7275258b",
   738 => x"38ad5195",
   739 => x"b12d7209",
   740 => x"81055372",
   741 => x"802eb538",
   742 => x"8754729c",
   743 => x"2a73842b",
   744 => x"54527180",
   745 => x"2e833881",
   746 => x"55897225",
   747 => x"8738b712",
   748 => x"5297b704",
   749 => x"b0125274",
   750 => x"802e8638",
   751 => x"715195b1",
   752 => x"2dff1454",
   753 => x"738025d2",
   754 => x"3897d104",
   755 => x"b05195b1",
   756 => x"2d800bb3",
   757 => x"e40c0294",
   758 => x"050d0402",
   759 => x"c0050d02",
   760 => x"80c40557",
   761 => x"80707870",
   762 => x"84055a08",
   763 => x"72415f5d",
   764 => x"587c7084",
   765 => x"055e085a",
   766 => x"805b7998",
   767 => x"2a7a882b",
   768 => x"5b567586",
   769 => x"38775f99",
   770 => x"d3047d80",
   771 => x"2e81a238",
   772 => x"805e7580",
   773 => x"e42e8a38",
   774 => x"7580f82e",
   775 => x"09810689",
   776 => x"38768418",
   777 => x"71085e58",
   778 => x"547580e4",
   779 => x"2e9f3875",
   780 => x"80e4268a",
   781 => x"387580e3",
   782 => x"2ebe3899",
   783 => x"83047580",
   784 => x"f32ea338",
   785 => x"7580f82e",
   786 => x"89389983",
   787 => x"048a5398",
   788 => x"d4049053",
   789 => x"b4c4527b",
   790 => x"5196fc2d",
   791 => x"b3e408b4",
   792 => x"c45a5599",
   793 => x"93047684",
   794 => x"18710870",
   795 => x"545b5854",
   796 => x"95d32d80",
   797 => x"55999304",
   798 => x"76841871",
   799 => x"08585854",
   800 => x"99be04a5",
   801 => x"5195b12d",
   802 => x"755195b1",
   803 => x"2d821858",
   804 => x"99c60474",
   805 => x"ff165654",
   806 => x"807425aa",
   807 => x"38787081",
   808 => x"055a80f5",
   809 => x"2d705256",
   810 => x"95b12d81",
   811 => x"18589993",
   812 => x"0475a52e",
   813 => x"09810686",
   814 => x"38815e99",
   815 => x"c6047551",
   816 => x"95b12d81",
   817 => x"1858811b",
   818 => x"5b837b25",
   819 => x"feac3875",
   820 => x"fe9f387e",
   821 => x"b3e40c02",
   822 => x"80c0050d",
   823 => x"0402ec05",
   824 => x"0d765574",
   825 => x"80f52d51",
   826 => x"70802e81",
   827 => x"f238b588",
   828 => x"08708280",
   829 => x"8029a9e0",
   830 => x"0805b584",
   831 => x"08115152",
   832 => x"52718f24",
   833 => x"de387470",
   834 => x"81055680",
   835 => x"f52d5271",
   836 => x"802e81cb",
   837 => x"3871882e",
   838 => x"0981069c",
   839 => x"38800bb5",
   840 => x"840825b8",
   841 => x"38ff1151",
   842 => x"a07181b7",
   843 => x"2db58408",
   844 => x"ff05b584",
   845 => x"0c9b8404",
   846 => x"718a2e09",
   847 => x"81069d38",
   848 => x"b5880881",
   849 => x"05b5880c",
   850 => x"800bb584",
   851 => x"0cb58808",
   852 => x"82808029",
   853 => x"a9e00805",
   854 => x"519b8404",
   855 => x"71717081",
   856 => x"055381b7",
   857 => x"2db58408",
   858 => x"8105b584",
   859 => x"0cb58408",
   860 => x"a02e0981",
   861 => x"068e3880",
   862 => x"0bb5840c",
   863 => x"b5880881",
   864 => x"05b5880c",
   865 => x"8f0bb588",
   866 => x"082580c7",
   867 => x"38a9e008",
   868 => x"82808011",
   869 => x"71535553",
   870 => x"81ff5273",
   871 => x"70840555",
   872 => x"08717084",
   873 => x"05530cff",
   874 => x"12527180",
   875 => x"25ed3888",
   876 => x"8013518f",
   877 => x"52807170",
   878 => x"8405530c",
   879 => x"ff125271",
   880 => x"8025f238",
   881 => x"800bb584",
   882 => x"0c8f0bb5",
   883 => x"880c9e80",
   884 => x"8013518f",
   885 => x"0bb58808",
   886 => x"25feab38",
   887 => x"99e30402",
   888 => x"94050d04",
   889 => x"02f4050d",
   890 => x"02930580",
   891 => x"f52d028c",
   892 => x"0581b72d",
   893 => x"80028405",
   894 => x"890581b7",
   895 => x"2d028c05",
   896 => x"fc055199",
   897 => x"dd2d810b",
   898 => x"b3e40c02",
   899 => x"8c050d04",
   900 => x"02fc050d",
   901 => x"725199dd",
   902 => x"2d800bb3",
   903 => x"e40c0284",
   904 => x"050d0402",
   905 => x"f8050da9",
   906 => x"e008528f",
   907 => x"fc518072",
   908 => x"70840554",
   909 => x"0cfc1151",
   910 => x"708025f2",
   911 => x"38028805",
   912 => x"0d0402fc",
   913 => x"050d7251",
   914 => x"80710c80",
   915 => x"0b84120c",
   916 => x"800b8812",
   917 => x"0c800b8c",
   918 => x"120c0284",
   919 => x"050d0402",
   920 => x"f0050d75",
   921 => x"70088412",
   922 => x"08535353",
   923 => x"ff547171",
   924 => x"2e9b3884",
   925 => x"13087084",
   926 => x"29149311",
   927 => x"80f52d84",
   928 => x"16088111",
   929 => x"87068418",
   930 => x"0c525651",
   931 => x"5173b3e4",
   932 => x"0c029005",
   933 => x"0d0402f4",
   934 => x"050d7470",
   935 => x"08841208",
   936 => x"53535370",
   937 => x"72248f38",
   938 => x"72088414",
   939 => x"08717131",
   940 => x"5252529d",
   941 => x"c3047208",
   942 => x"84140871",
   943 => x"71318805",
   944 => x"52525271",
   945 => x"b3e40c02",
   946 => x"8c050d04",
   947 => x"02f8050d",
   948 => x"a2b02da2",
   949 => x"a32de008",
   950 => x"708b2a70",
   951 => x"81065152",
   952 => x"5270802e",
   953 => x"9d38b9ec",
   954 => x"08708429",
   955 => x"b9fc0573",
   956 => x"81ff0671",
   957 => x"0c5151b9",
   958 => x"ec088111",
   959 => x"8706b9ec",
   960 => x"0c51718a",
   961 => x"2a708106",
   962 => x"51517080",
   963 => x"2ea838b9",
   964 => x"f408b9f8",
   965 => x"08525271",
   966 => x"712e9b38",
   967 => x"b9f40870",
   968 => x"8429ba9c",
   969 => x"057008e0",
   970 => x"0c5151b9",
   971 => x"f4088111",
   972 => x"8706b9f4",
   973 => x"0c51a2aa",
   974 => x"2d028805",
   975 => x"0d0402f4",
   976 => x"050d7453",
   977 => x"8c130881",
   978 => x"11870688",
   979 => x"15085451",
   980 => x"5171712e",
   981 => x"ef38a2b0",
   982 => x"2d8c1308",
   983 => x"70842914",
   984 => x"77b0120c",
   985 => x"51518c13",
   986 => x"08811187",
   987 => x"068c150c",
   988 => x"519dcc2d",
   989 => x"a2aa2d02",
   990 => x"8c050d04",
   991 => x"02fc050d",
   992 => x"b9ec519c",
   993 => x"c22d9dcc",
   994 => x"51a29f2d",
   995 => x"a1d72d02",
   996 => x"84050d04",
   997 => x"02e4050d",
   998 => x"8057a1a2",
   999 => x"04b3e408",
  1000 => x"81f02e09",
  1001 => x"81068938",
  1002 => x"810bb594",
  1003 => x"0ca1a204",
  1004 => x"b3e40881",
  1005 => x"e02e0981",
  1006 => x"06893881",
  1007 => x"0bb5980c",
  1008 => x"a1a204b3",
  1009 => x"e40854b5",
  1010 => x"9808802e",
  1011 => x"8838b3e4",
  1012 => x"08818005",
  1013 => x"54b59408",
  1014 => x"819c3883",
  1015 => x"0ba9e415",
  1016 => x"81b72d74",
  1017 => x"80ff24b1",
  1018 => x"38b59008",
  1019 => x"822a7081",
  1020 => x"06b58c08",
  1021 => x"70872b81",
  1022 => x"80077811",
  1023 => x"822b5156",
  1024 => x"58515473",
  1025 => x"8b387581",
  1026 => x"80291570",
  1027 => x"822b5153",
  1028 => x"abe41308",
  1029 => x"537281b6",
  1030 => x"38800bb5",
  1031 => x"980c7480",
  1032 => x"d92e80c7",
  1033 => x"387480d9",
  1034 => x"248f3874",
  1035 => x"922ebc38",
  1036 => x"7480d82e",
  1037 => x"9338a19d",
  1038 => x"047480f7",
  1039 => x"2ea03874",
  1040 => x"80fe2e8f",
  1041 => x"38a19d04",
  1042 => x"b5900884",
  1043 => x"32b5900c",
  1044 => x"a0e604b5",
  1045 => x"90088132",
  1046 => x"b5900ca0",
  1047 => x"e604b590",
  1048 => x"088232b5",
  1049 => x"900c8157",
  1050 => x"a19d04b5",
  1051 => x"8c088107",
  1052 => x"b58c0ca1",
  1053 => x"9d04a9e4",
  1054 => x"1480f52d",
  1055 => x"81fe0653",
  1056 => x"72a9e415",
  1057 => x"81b72d74",
  1058 => x"922e8a38",
  1059 => x"7480d92e",
  1060 => x"09810689",
  1061 => x"38b58c08",
  1062 => x"fe06b58c",
  1063 => x"0c800bb5",
  1064 => x"940cb9ec",
  1065 => x"519cdf2d",
  1066 => x"b3e40855",
  1067 => x"b3e408ff",
  1068 => x"24fdea38",
  1069 => x"76802e94",
  1070 => x"3881ed52",
  1071 => x"b9ec519e",
  1072 => x"be2db590",
  1073 => x"0852b9ec",
  1074 => x"519ebe2d",
  1075 => x"805372b3",
  1076 => x"e40c029c",
  1077 => x"050d0402",
  1078 => x"fc050d80",
  1079 => x"51800ba9",
  1080 => x"e41281b7",
  1081 => x"2d811151",
  1082 => x"81ff7125",
  1083 => x"f0380284",
  1084 => x"050d0402",
  1085 => x"f4050d74",
  1086 => x"51a2b02d",
  1087 => x"a9e41180",
  1088 => x"f52d7081",
  1089 => x"ff0671fd",
  1090 => x"06525452",
  1091 => x"71a9e412",
  1092 => x"81b72da2",
  1093 => x"aa2d72b3",
  1094 => x"e40c028c",
  1095 => x"050d0471",
  1096 => x"980c04ff",
  1097 => x"b008b3e4",
  1098 => x"0c04810b",
  1099 => x"ffb00c04",
  1100 => x"800bffb0",
  1101 => x"0c0402e8",
  1102 => x"050d7878",
  1103 => x"71545753",
  1104 => x"72802584",
  1105 => x"38831352",
  1106 => x"71822cff",
  1107 => x"055372ff",
  1108 => x"2e80c038",
  1109 => x"75708405",
  1110 => x"57085487",
  1111 => x"55739c2a",
  1112 => x"b00552b9",
  1113 => x"72278438",
  1114 => x"87125271",
  1115 => x"5195b12d",
  1116 => x"73842bff",
  1117 => x"16565474",
  1118 => x"8025e238",
  1119 => x"a05195b1",
  1120 => x"2d728706",
  1121 => x"52718638",
  1122 => x"8a5195b1",
  1123 => x"2dff1353",
  1124 => x"a2ce048a",
  1125 => x"5195b12d",
  1126 => x"0298050d",
  1127 => x"04b3f008",
  1128 => x"02b3f00c",
  1129 => x"ff3d0d80",
  1130 => x"0bb3f008",
  1131 => x"fc050cb3",
  1132 => x"f0088805",
  1133 => x"088106ff",
  1134 => x"11700970",
  1135 => x"b3f0088c",
  1136 => x"050806b3",
  1137 => x"f008fc05",
  1138 => x"0811b3f0",
  1139 => x"08fc050c",
  1140 => x"b3f00888",
  1141 => x"0508812a",
  1142 => x"b3f00888",
  1143 => x"050cb3f0",
  1144 => x"088c0508",
  1145 => x"10b3f008",
  1146 => x"8c050c51",
  1147 => x"515151b3",
  1148 => x"f0088805",
  1149 => x"08802e84",
  1150 => x"38ffb439",
  1151 => x"b3f008fc",
  1152 => x"050870b3",
  1153 => x"e40c5183",
  1154 => x"3d0db3f0",
  1155 => x"0c040000",
  1156 => x"00ffffff",
  1157 => x"ff00ffff",
  1158 => x"ffff00ff",
  1159 => x"ffffff00",
  1160 => x"496e6974",
  1161 => x"69616c69",
  1162 => x"73696e67",
  1163 => x"2050532f",
  1164 => x"3220696e",
  1165 => x"74657266",
  1166 => x"6163652e",
  1167 => x"2e2e0a00",
  1168 => x"496e6974",
  1169 => x"69616c69",
  1170 => x"7a696e67",
  1171 => x"20534420",
  1172 => x"63617264",
  1173 => x"0a000000",
  1174 => x"48756e74",
  1175 => x"696e6720",
  1176 => x"666f7220",
  1177 => x"70617274",
  1178 => x"6974696f",
  1179 => x"6e0a0000",
  1180 => x"42494f53",
  1181 => x"5f4d3250",
  1182 => x"524f4d00",
  1183 => x"4f70656e",
  1184 => x"65642066",
  1185 => x"696c652c",
  1186 => x"206c6f61",
  1187 => x"64696e67",
  1188 => x"2e2e2e0a",
  1189 => x"00000000",
  1190 => x"52656164",
  1191 => x"20626c6f",
  1192 => x"636b2066",
  1193 => x"61696c65",
  1194 => x"640a0000",
  1195 => x"4c6f6164",
  1196 => x"696e6720",
  1197 => x"42494f53",
  1198 => x"20666169",
  1199 => x"6c65640a",
  1200 => x"00000000",
  1201 => x"52656164",
  1202 => x"696e6720",
  1203 => x"4d42520a",
  1204 => x"00000000",
  1205 => x"52656164",
  1206 => x"206f6620",
  1207 => x"4d425220",
  1208 => x"6661696c",
  1209 => x"65640a00",
  1210 => x"4d425220",
  1211 => x"73756363",
  1212 => x"65737366",
  1213 => x"756c6c79",
  1214 => x"20726561",
  1215 => x"640a0000",
  1216 => x"46415431",
  1217 => x"36202020",
  1218 => x"00000000",
  1219 => x"46415433",
  1220 => x"32202020",
  1221 => x"00000000",
  1222 => x"50617274",
  1223 => x"6974696f",
  1224 => x"6e636f75",
  1225 => x"6e742025",
  1226 => x"640a0000",
  1227 => x"4e6f2070",
  1228 => x"61727469",
  1229 => x"74696f6e",
  1230 => x"20736967",
  1231 => x"6e617475",
  1232 => x"72652066",
  1233 => x"6f756e64",
  1234 => x"0a000000",
  1235 => x"52656164",
  1236 => x"696e6720",
  1237 => x"626f6f74",
  1238 => x"20736563",
  1239 => x"746f7220",
  1240 => x"25640a00",
  1241 => x"52656164",
  1242 => x"20626f6f",
  1243 => x"74207365",
  1244 => x"63746f72",
  1245 => x"2066726f",
  1246 => x"6d206669",
  1247 => x"72737420",
  1248 => x"70617274",
  1249 => x"6974696f",
  1250 => x"6e0a0000",
  1251 => x"48756e74",
  1252 => x"696e6720",
  1253 => x"666f7220",
  1254 => x"66696c65",
  1255 => x"73797374",
  1256 => x"656d0a00",
  1257 => x"556e7375",
  1258 => x"70706f72",
  1259 => x"74656420",
  1260 => x"70617274",
  1261 => x"6974696f",
  1262 => x"6e207479",
  1263 => x"7065210d",
  1264 => x"00000000",
  1265 => x"436c7573",
  1266 => x"74657220",
  1267 => x"73697a65",
  1268 => x"3a202564",
  1269 => x"2c20436c",
  1270 => x"75737465",
  1271 => x"72206d61",
  1272 => x"736b2c20",
  1273 => x"25640a00",
  1274 => x"47657443",
  1275 => x"6c757374",
  1276 => x"65722072",
  1277 => x"65616469",
  1278 => x"6e672073",
  1279 => x"6563746f",
  1280 => x"72202564",
  1281 => x"0a000000",
  1282 => x"52656164",
  1283 => x"696e6720",
  1284 => x"64697265",
  1285 => x"63746f72",
  1286 => x"79207365",
  1287 => x"63746f72",
  1288 => x"2025640a",
  1289 => x"00000000",
  1290 => x"47657446",
  1291 => x"41544c69",
  1292 => x"6e6b2072",
  1293 => x"65747572",
  1294 => x"6e656420",
  1295 => x"25640a00",
  1296 => x"436d645f",
  1297 => x"696e6974",
  1298 => x"0a000000",
  1299 => x"636d645f",
  1300 => x"434d4438",
  1301 => x"20726573",
  1302 => x"706f6e73",
  1303 => x"653a2025",
  1304 => x"640a0000",
  1305 => x"434d4438",
  1306 => x"5f342072",
  1307 => x"6573706f",
  1308 => x"6e73653a",
  1309 => x"2025640a",
  1310 => x"00000000",
  1311 => x"53444843",
  1312 => x"20496e69",
  1313 => x"7469616c",
  1314 => x"697a6174",
  1315 => x"696f6e20",
  1316 => x"6572726f",
  1317 => x"72210a00",
  1318 => x"434d4435",
  1319 => x"38202564",
  1320 => x"0a202000",
  1321 => x"434d4435",
  1322 => x"385f3220",
  1323 => x"25640a20",
  1324 => x"20000000",
  1325 => x"53504920",
  1326 => x"496e6974",
  1327 => x"28290a00",
  1328 => x"52656164",
  1329 => x"20636f6d",
  1330 => x"6d616e64",
  1331 => x"20666169",
  1332 => x"6c656420",
  1333 => x"61742025",
  1334 => x"64202825",
  1335 => x"64290a00",
  1336 => x"ffffe000",
  1337 => x"00000000",
  1338 => x"00000000",
  1339 => x"00000000",
  1340 => x"00000000",
  1341 => x"00000000",
  1342 => x"00000000",
  1343 => x"00000000",
  1344 => x"00000000",
  1345 => x"00000000",
  1346 => x"00000000",
  1347 => x"00000000",
  1348 => x"00000000",
  1349 => x"00000000",
  1350 => x"00000000",
  1351 => x"00000000",
  1352 => x"00000000",
  1353 => x"00000000",
  1354 => x"00000000",
  1355 => x"00000000",
  1356 => x"00000000",
  1357 => x"00000000",
  1358 => x"00000000",
  1359 => x"00000000",
  1360 => x"00000000",
  1361 => x"00000000",
  1362 => x"00000000",
  1363 => x"00000000",
  1364 => x"00000000",
  1365 => x"00000000",
  1366 => x"00000000",
  1367 => x"00000000",
  1368 => x"00000000",
  1369 => x"00000000",
  1370 => x"00000000",
  1371 => x"00000000",
  1372 => x"00000000",
  1373 => x"00000000",
  1374 => x"00000000",
  1375 => x"00000000",
  1376 => x"00000000",
  1377 => x"00000000",
  1378 => x"00000000",
  1379 => x"00000000",
  1380 => x"00000000",
  1381 => x"00000000",
  1382 => x"00000000",
  1383 => x"00000000",
  1384 => x"00000000",
  1385 => x"00000000",
  1386 => x"00000000",
  1387 => x"00000000",
  1388 => x"00000000",
  1389 => x"00000000",
  1390 => x"00000000",
  1391 => x"00000000",
  1392 => x"00000000",
  1393 => x"00000000",
  1394 => x"00000000",
  1395 => x"00000000",
  1396 => x"00000000",
  1397 => x"00000000",
  1398 => x"00000000",
  1399 => x"00000000",
  1400 => x"00000000",
  1401 => x"00000000",
  1402 => x"00000000",
  1403 => x"00000000",
  1404 => x"00000000",
  1405 => x"00000000",
  1406 => x"00000000",
  1407 => x"00000000",
  1408 => x"00000000",
  1409 => x"00000000",
  1410 => x"00000000",
  1411 => x"00000000",
  1412 => x"00000000",
  1413 => x"00000000",
  1414 => x"00000009",
  1415 => x"00000000",
  1416 => x"00000000",
  1417 => x"00000000",
  1418 => x"00000000",
  1419 => x"00000000",
  1420 => x"00000000",
  1421 => x"00000000",
  1422 => x"00000071",
  1423 => x"00000031",
  1424 => x"00000000",
  1425 => x"00000000",
  1426 => x"00000000",
  1427 => x"0000007a",
  1428 => x"00000073",
  1429 => x"00000061",
  1430 => x"00000077",
  1431 => x"00000032",
  1432 => x"00000000",
  1433 => x"00000000",
  1434 => x"00000063",
  1435 => x"00000078",
  1436 => x"00000064",
  1437 => x"00000065",
  1438 => x"00000034",
  1439 => x"00000033",
  1440 => x"00000000",
  1441 => x"00000000",
  1442 => x"00000020",
  1443 => x"00000076",
  1444 => x"00000066",
  1445 => x"00000074",
  1446 => x"00000072",
  1447 => x"00000035",
  1448 => x"00000000",
  1449 => x"00000000",
  1450 => x"0000006e",
  1451 => x"00000062",
  1452 => x"00000068",
  1453 => x"00000067",
  1454 => x"00000079",
  1455 => x"00000036",
  1456 => x"00000000",
  1457 => x"00000000",
  1458 => x"00000000",
  1459 => x"0000006d",
  1460 => x"0000006a",
  1461 => x"00000075",
  1462 => x"00000037",
  1463 => x"00000038",
  1464 => x"00000000",
  1465 => x"00000000",
  1466 => x"0000002c",
  1467 => x"0000006b",
  1468 => x"00000069",
  1469 => x"0000006f",
  1470 => x"00000030",
  1471 => x"00000039",
  1472 => x"00000000",
  1473 => x"00000000",
  1474 => x"0000002e",
  1475 => x"0000002f",
  1476 => x"0000006c",
  1477 => x"0000003b",
  1478 => x"00000070",
  1479 => x"0000002d",
  1480 => x"00000000",
  1481 => x"00000000",
  1482 => x"00000000",
  1483 => x"00000027",
  1484 => x"00000000",
  1485 => x"0000005b",
  1486 => x"0000003d",
  1487 => x"00000000",
  1488 => x"00000000",
  1489 => x"00000000",
  1490 => x"00000000",
  1491 => x"0000000a",
  1492 => x"0000005d",
  1493 => x"00000000",
  1494 => x"00000023",
  1495 => x"00000000",
  1496 => x"00000000",
  1497 => x"00000000",
  1498 => x"00000000",
  1499 => x"00000000",
  1500 => x"00000000",
  1501 => x"00000000",
  1502 => x"00000000",
  1503 => x"00000008",
  1504 => x"00000000",
  1505 => x"00000000",
  1506 => x"00000031",
  1507 => x"00000000",
  1508 => x"00000034",
  1509 => x"00000037",
  1510 => x"00000000",
  1511 => x"00000000",
  1512 => x"00000000",
  1513 => x"00000030",
  1514 => x"0000002e",
  1515 => x"00000032",
  1516 => x"00000035",
  1517 => x"00000036",
  1518 => x"00000038",
  1519 => x"0000001b",
  1520 => x"00000000",
  1521 => x"00000000",
  1522 => x"0000002b",
  1523 => x"00000033",
  1524 => x"00000000",
  1525 => x"0000002a",
  1526 => x"00000039",
  1527 => x"00000000",
  1528 => x"00000000",
  1529 => x"00000000",
  1530 => x"00000000",
  1531 => x"00000000",
  1532 => x"00000000",
  1533 => x"00000000",
  1534 => x"00000000",
  1535 => x"00000000",
  1536 => x"00000000",
  1537 => x"00000000",
  1538 => x"00000000",
  1539 => x"00000000",
  1540 => x"00000000",
  1541 => x"00000000",
  1542 => x"00000008",
  1543 => x"00000000",
  1544 => x"00000000",
  1545 => x"00000000",
  1546 => x"00000000",
  1547 => x"00000000",
  1548 => x"00000000",
  1549 => x"00000000",
  1550 => x"00000051",
  1551 => x"00000021",
  1552 => x"00000000",
  1553 => x"00000000",
  1554 => x"00000000",
  1555 => x"0000005a",
  1556 => x"00000053",
  1557 => x"00000041",
  1558 => x"00000057",
  1559 => x"00000022",
  1560 => x"00000000",
  1561 => x"00000000",
  1562 => x"00000043",
  1563 => x"00000058",
  1564 => x"00000044",
  1565 => x"00000045",
  1566 => x"00000024",
  1567 => x"000000a3",
  1568 => x"00000000",
  1569 => x"00000000",
  1570 => x"00000020",
  1571 => x"00000056",
  1572 => x"00000046",
  1573 => x"00000054",
  1574 => x"00000052",
  1575 => x"00000025",
  1576 => x"00000000",
  1577 => x"00000000",
  1578 => x"0000004e",
  1579 => x"00000042",
  1580 => x"00000048",
  1581 => x"00000047",
  1582 => x"00000059",
  1583 => x"0000005e",
  1584 => x"00000000",
  1585 => x"00000000",
  1586 => x"00000000",
  1587 => x"0000004d",
  1588 => x"0000004a",
  1589 => x"00000055",
  1590 => x"00000026",
  1591 => x"0000002a",
  1592 => x"00000000",
  1593 => x"00000000",
  1594 => x"0000003c",
  1595 => x"0000004b",
  1596 => x"00000049",
  1597 => x"0000004f",
  1598 => x"00000029",
  1599 => x"00000028",
  1600 => x"00000000",
  1601 => x"00000000",
  1602 => x"0000003e",
  1603 => x"0000003f",
  1604 => x"0000004c",
  1605 => x"0000003a",
  1606 => x"00000050",
  1607 => x"0000005f",
  1608 => x"00000000",
  1609 => x"00000000",
  1610 => x"00000000",
  1611 => x"0000003f",
  1612 => x"00000000",
  1613 => x"0000007b",
  1614 => x"0000002b",
  1615 => x"00000000",
  1616 => x"00000000",
  1617 => x"00000000",
  1618 => x"00000000",
  1619 => x"0000000a",
  1620 => x"0000007d",
  1621 => x"00000000",
  1622 => x"0000007e",
  1623 => x"00000000",
  1624 => x"00000000",
  1625 => x"00000000",
  1626 => x"00000000",
  1627 => x"00000000",
  1628 => x"00000000",
  1629 => x"00000000",
  1630 => x"00000000",
  1631 => x"00000009",
  1632 => x"00000000",
  1633 => x"00000000",
  1634 => x"00000031",
  1635 => x"00000000",
  1636 => x"00000034",
  1637 => x"00000037",
  1638 => x"00000000",
  1639 => x"00000000",
  1640 => x"00000000",
  1641 => x"00000030",
  1642 => x"0000002e",
  1643 => x"00000032",
  1644 => x"00000035",
  1645 => x"00000036",
  1646 => x"00000038",
  1647 => x"0000001b",
  1648 => x"00000000",
  1649 => x"00000000",
  1650 => x"0000002b",
  1651 => x"00000033",
  1652 => x"00000000",
  1653 => x"0000002a",
  1654 => x"00000039",
  1655 => x"00000000",
  1656 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

