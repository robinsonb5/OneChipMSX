-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b0bae",
     9 => x"e0080b0b",
    10 => x"0baee408",
    11 => x"0b0b0bae",
    12 => x"e8080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"aee80c0b",
    16 => x"0b0baee4",
    17 => x"0c0b0b0b",
    18 => x"aee00c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0ba5b0",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"aee070b4",
    57 => x"bc278b38",
    58 => x"80717084",
    59 => x"05530c81",
    60 => x"e2048c51",
    61 => x"86b30402",
    62 => x"fc050df8",
    63 => x"80518f0b",
    64 => x"aef00c9f",
    65 => x"0baef40c",
    66 => x"a0717081",
    67 => x"055334ae",
    68 => x"f408ff05",
    69 => x"aef40cae",
    70 => x"f4088025",
    71 => x"eb38aef0",
    72 => x"08ff05ae",
    73 => x"f00caef0",
    74 => x"088025d7",
    75 => x"38028405",
    76 => x"0d0402f0",
    77 => x"050df880",
    78 => x"53f8a054",
    79 => x"83bf5273",
    80 => x"70810555",
    81 => x"33517073",
    82 => x"70810555",
    83 => x"34ff1252",
    84 => x"718025eb",
    85 => x"38fbc053",
    86 => x"9f52a073",
    87 => x"70810555",
    88 => x"34ff1252",
    89 => x"718025f2",
    90 => x"38029005",
    91 => x"0d0402f4",
    92 => x"050d7453",
    93 => x"8e0baef0",
    94 => x"08258f38",
    95 => x"82b22dae",
    96 => x"f008ff05",
    97 => x"aef00c82",
    98 => x"f404aef0",
    99 => x"08aef408",
   100 => x"5351728a",
   101 => x"2e098106",
   102 => x"b7387151",
   103 => x"719f24a0",
   104 => x"38aef008",
   105 => x"a02911f8",
   106 => x"80115151",
   107 => x"a07134ae",
   108 => x"f4088105",
   109 => x"aef40cae",
   110 => x"f408519f",
   111 => x"7125e238",
   112 => x"800baef4",
   113 => x"0caef008",
   114 => x"8105aef0",
   115 => x"0c83e404",
   116 => x"70a02912",
   117 => x"f8801151",
   118 => x"51727134",
   119 => x"aef40881",
   120 => x"05aef40c",
   121 => x"aef408a0",
   122 => x"2e098106",
   123 => x"8e38800b",
   124 => x"aef40cae",
   125 => x"f0088105",
   126 => x"aef00c02",
   127 => x"8c050d04",
   128 => x"02e8050d",
   129 => x"77795656",
   130 => x"880bfc16",
   131 => x"77712c8f",
   132 => x"06545254",
   133 => x"80537272",
   134 => x"25953871",
   135 => x"53fbe014",
   136 => x"51877134",
   137 => x"8114ff14",
   138 => x"545472f1",
   139 => x"387153f9",
   140 => x"1576712c",
   141 => x"87065351",
   142 => x"71802e8b",
   143 => x"38fbe014",
   144 => x"51717134",
   145 => x"81145472",
   146 => x"8e249538",
   147 => x"8f733153",
   148 => x"fbe01451",
   149 => x"a0713481",
   150 => x"14ff1454",
   151 => x"5472f138",
   152 => x"0298050d",
   153 => x"0402ec05",
   154 => x"0d800bae",
   155 => x"fc0cf68c",
   156 => x"08f69008",
   157 => x"71882c57",
   158 => x"5481ff06",
   159 => x"52747225",
   160 => x"88387155",
   161 => x"820baefc",
   162 => x"0c72882c",
   163 => x"7381ff06",
   164 => x"54547373",
   165 => x"258b3872",
   166 => x"aefc0884",
   167 => x"07aefc0c",
   168 => x"54aef808",
   169 => x"82055182",
   170 => x"0baef80c",
   171 => x"830bf688",
   172 => x"0c74712b",
   173 => x"fecc0570",
   174 => x"9f2a1170",
   175 => x"812c7688",
   176 => x"29ff9405",
   177 => x"70812cae",
   178 => x"fc085257",
   179 => x"52545151",
   180 => x"76802e85",
   181 => x"38708107",
   182 => x"5170f694",
   183 => x"0c710981",
   184 => x"05f6800c",
   185 => x"72098105",
   186 => x"f6840c02",
   187 => x"94050d04",
   188 => x"02f4050d",
   189 => x"74537270",
   190 => x"81055480",
   191 => x"f52d5271",
   192 => x"802e8938",
   193 => x"715182ee",
   194 => x"2d85f604",
   195 => x"028c050d",
   196 => x"040402f8",
   197 => x"050d9fb5",
   198 => x"2d80da51",
   199 => x"a0ec2dae",
   200 => x"e008812a",
   201 => x"70810651",
   202 => x"5271802e",
   203 => x"e9380288",
   204 => x"050d0402",
   205 => x"d4050d81",
   206 => x"0bfec40c",
   207 => x"b90bfec0",
   208 => x"0c840bfe",
   209 => x"c40c9f9d",
   210 => x"2da1b02d",
   211 => x"9f822d9f",
   212 => x"822d81f7",
   213 => x"2d815184",
   214 => x"e52d9f82",
   215 => x"2d9f822d",
   216 => x"815184e5",
   217 => x"2da89451",
   218 => x"85f02d97",
   219 => x"bd2daee0",
   220 => x"08802e82",
   221 => x"ad3889f0",
   222 => x"2daee008",
   223 => x"53aee008",
   224 => x"802e82a5",
   225 => x"3899f92d",
   226 => x"aee00880",
   227 => x"2e8738a8",
   228 => x"ac5187a2",
   229 => x"0493882d",
   230 => x"aee00880",
   231 => x"2e8a38a8",
   232 => x"ec5185f0",
   233 => x"2d86922d",
   234 => x"a9b45185",
   235 => x"f02da9cc",
   236 => x"52af8051",
   237 => x"908c2dae",
   238 => x"e00881ff",
   239 => x"0653729d",
   240 => x"38a9d851",
   241 => x"85f02da9",
   242 => x"f052af80",
   243 => x"51908c2d",
   244 => x"aee00881",
   245 => x"ff065372",
   246 => x"802e81c0",
   247 => x"38a9fc51",
   248 => x"85f02daf",
   249 => x"84085780",
   250 => x"77595a76",
   251 => x"7a2e8b38",
   252 => x"811a7881",
   253 => x"2a595a77",
   254 => x"f738f71a",
   255 => x"5a807725",
   256 => x"80fe3879",
   257 => x"52775184",
   258 => x"802daf8c",
   259 => x"52af8051",
   260 => x"92d12dae",
   261 => x"e00881ff",
   262 => x"06af8c5c",
   263 => x"53805972",
   264 => x"792e0981",
   265 => x"06b13888",
   266 => x"ea047a70",
   267 => x"84055c08",
   268 => x"7081ff06",
   269 => x"71882c70",
   270 => x"81ff0673",
   271 => x"902c7081",
   272 => x"ff067598",
   273 => x"2afec80c",
   274 => x"fec80c58",
   275 => x"fec80c57",
   276 => x"fec80c84",
   277 => x"1a5a5376",
   278 => x"53848077",
   279 => x"25843884",
   280 => x"80537279",
   281 => x"24c43888",
   282 => x"f004aa98",
   283 => x"519a802d",
   284 => x"af805192",
   285 => x"a42dfc80",
   286 => x"17811959",
   287 => x"5787fd04",
   288 => x"820bfec4",
   289 => x"0c805184",
   290 => x"e52d0b0b",
   291 => x"0bacc451",
   292 => x"a2d52d9f",
   293 => x"b52da2e5",
   294 => x"2d899304",
   295 => x"aaac519a",
   296 => x"802d820b",
   297 => x"fec40c80",
   298 => x"5372aee0",
   299 => x"0c02ac05",
   300 => x"0d0402e8",
   301 => x"050d7779",
   302 => x"7b585555",
   303 => x"80537276",
   304 => x"25a33874",
   305 => x"70810556",
   306 => x"80f52d74",
   307 => x"70810556",
   308 => x"80f52d52",
   309 => x"5271712e",
   310 => x"86388151",
   311 => x"89e70481",
   312 => x"135389be",
   313 => x"04805170",
   314 => x"aee00c02",
   315 => x"98050d04",
   316 => x"02d8050d",
   317 => x"800bb394",
   318 => x"0caf8c52",
   319 => x"805198d6",
   320 => x"2daee008",
   321 => x"54aee008",
   322 => x"8c38aac4",
   323 => x"5185f02d",
   324 => x"73558f95",
   325 => x"04805681",
   326 => x"0bb3b80c",
   327 => x"8853aad8",
   328 => x"52afc251",
   329 => x"89b22dae",
   330 => x"e008762e",
   331 => x"09810687",
   332 => x"38aee008",
   333 => x"b3b80c88",
   334 => x"53aae452",
   335 => x"afde5189",
   336 => x"b22daee0",
   337 => x"088738ae",
   338 => x"e008b3b8",
   339 => x"0cb3b808",
   340 => x"52aaf051",
   341 => x"9bf32db3",
   342 => x"b808802e",
   343 => x"80f638b2",
   344 => x"d20b80f5",
   345 => x"2db2d30b",
   346 => x"80f52d71",
   347 => x"982b7190",
   348 => x"2b07b2d4",
   349 => x"0b80f52d",
   350 => x"70882b72",
   351 => x"07b2d50b",
   352 => x"80f52d71",
   353 => x"07b38a0b",
   354 => x"80f52db3",
   355 => x"8b0b80f5",
   356 => x"2d71882b",
   357 => x"07535f54",
   358 => x"525a5657",
   359 => x"557381ab",
   360 => x"aa2e0981",
   361 => x"068d3875",
   362 => x"519ac82d",
   363 => x"aee00856",
   364 => x"8bc00473",
   365 => x"82d4d52e",
   366 => x"8738ab88",
   367 => x"518c8104",
   368 => x"af8c5275",
   369 => x"5198d62d",
   370 => x"aee00855",
   371 => x"aee00880",
   372 => x"2e83c238",
   373 => x"8853aae4",
   374 => x"52afde51",
   375 => x"89b22dae",
   376 => x"e0088938",
   377 => x"810bb394",
   378 => x"0c8c8704",
   379 => x"8853aad8",
   380 => x"52afc251",
   381 => x"89b22dae",
   382 => x"e008802e",
   383 => x"8a38aba8",
   384 => x"5185f02d",
   385 => x"8ce104b3",
   386 => x"8a0b80f5",
   387 => x"2d547380",
   388 => x"d52e0981",
   389 => x"0680ca38",
   390 => x"b38b0b80",
   391 => x"f52d5473",
   392 => x"81aa2e09",
   393 => x"8106ba38",
   394 => x"800baf8c",
   395 => x"0b80f52d",
   396 => x"56547481",
   397 => x"e92e8338",
   398 => x"81547481",
   399 => x"eb2e8c38",
   400 => x"80557375",
   401 => x"2e098106",
   402 => x"82cb38af",
   403 => x"970b80f5",
   404 => x"2d55748d",
   405 => x"38af980b",
   406 => x"80f52d54",
   407 => x"73822e86",
   408 => x"3880558f",
   409 => x"9504af99",
   410 => x"0b80f52d",
   411 => x"70b38c0c",
   412 => x"ff05b390",
   413 => x"0caf9a0b",
   414 => x"80f52daf",
   415 => x"9b0b80f5",
   416 => x"2d587605",
   417 => x"77828029",
   418 => x"0570b398",
   419 => x"0caf9c0b",
   420 => x"80f52d70",
   421 => x"b3ac0cb3",
   422 => x"94085957",
   423 => x"5876802e",
   424 => x"81a33888",
   425 => x"53aae452",
   426 => x"afde5189",
   427 => x"b22daee0",
   428 => x"0881e238",
   429 => x"b38c0870",
   430 => x"842bb3b0",
   431 => x"0c70b3a8",
   432 => x"0cafb10b",
   433 => x"80f52daf",
   434 => x"b00b80f5",
   435 => x"2d718280",
   436 => x"2905afb2",
   437 => x"0b80f52d",
   438 => x"70848080",
   439 => x"2912afb3",
   440 => x"0b80f52d",
   441 => x"7081800a",
   442 => x"291270b3",
   443 => x"b40cb3ac",
   444 => x"087129b3",
   445 => x"98080570",
   446 => x"b39c0caf",
   447 => x"b90b80f5",
   448 => x"2dafb80b",
   449 => x"80f52d71",
   450 => x"82802905",
   451 => x"afba0b80",
   452 => x"f52d7084",
   453 => x"80802912",
   454 => x"afbb0b80",
   455 => x"f52d7098",
   456 => x"2b81f00a",
   457 => x"06720570",
   458 => x"b3a00cfe",
   459 => x"117e2977",
   460 => x"05b3a40c",
   461 => x"52595243",
   462 => x"545e5152",
   463 => x"59525d57",
   464 => x"59578f93",
   465 => x"04af9e0b",
   466 => x"80f52daf",
   467 => x"9d0b80f5",
   468 => x"2d718280",
   469 => x"290570b3",
   470 => x"b00c70a0",
   471 => x"2983ff05",
   472 => x"70892a70",
   473 => x"b3a80caf",
   474 => x"a30b80f5",
   475 => x"2dafa20b",
   476 => x"80f52d71",
   477 => x"82802905",
   478 => x"70b3b40c",
   479 => x"7b71291e",
   480 => x"70b3a40c",
   481 => x"7db3a00c",
   482 => x"7305b39c",
   483 => x"0c555e51",
   484 => x"51555581",
   485 => x"5574aee0",
   486 => x"0c02a805",
   487 => x"0d0402ec",
   488 => x"050d7670",
   489 => x"872c7180",
   490 => x"ff065556",
   491 => x"54b39408",
   492 => x"8a387388",
   493 => x"2c7481ff",
   494 => x"065455af",
   495 => x"8c52b398",
   496 => x"08155198",
   497 => x"d62daee0",
   498 => x"0854aee0",
   499 => x"08802eb3",
   500 => x"38b39408",
   501 => x"802e9838",
   502 => x"728429af",
   503 => x"8c057008",
   504 => x"52539ac8",
   505 => x"2daee008",
   506 => x"f00a0653",
   507 => x"90810472",
   508 => x"10af8c05",
   509 => x"7080e02d",
   510 => x"52539af8",
   511 => x"2daee008",
   512 => x"53725473",
   513 => x"aee00c02",
   514 => x"94050d04",
   515 => x"02c8050d",
   516 => x"7f615f5b",
   517 => x"800bb3a0",
   518 => x"08b3a408",
   519 => x"595d56b3",
   520 => x"9408762e",
   521 => x"8a38b38c",
   522 => x"08842b58",
   523 => x"90b504b3",
   524 => x"a808842b",
   525 => x"58805978",
   526 => x"782781a9",
   527 => x"38788f06",
   528 => x"a0175754",
   529 => x"738f38af",
   530 => x"8c527651",
   531 => x"81175798",
   532 => x"d62daf8c",
   533 => x"56807680",
   534 => x"f52d5654",
   535 => x"74742e83",
   536 => x"38815474",
   537 => x"81e52e80",
   538 => x"f6388170",
   539 => x"7506555d",
   540 => x"73802e80",
   541 => x"ea388b16",
   542 => x"80f52d98",
   543 => x"065a7980",
   544 => x"de388b53",
   545 => x"7d527551",
   546 => x"89b22dae",
   547 => x"e00880cf",
   548 => x"389c1608",
   549 => x"519ac82d",
   550 => x"aee00884",
   551 => x"1c0c9a16",
   552 => x"80e02d51",
   553 => x"9af82dae",
   554 => x"e008aee0",
   555 => x"08881d0c",
   556 => x"aee00855",
   557 => x"55b39408",
   558 => x"802e9838",
   559 => x"941680e0",
   560 => x"2d519af8",
   561 => x"2daee008",
   562 => x"902b83ff",
   563 => x"f00a0670",
   564 => x"16515473",
   565 => x"881c0c79",
   566 => x"7b0c7c54",
   567 => x"929b0481",
   568 => x"195990b7",
   569 => x"04b39408",
   570 => x"802eae38",
   571 => x"7b518f9e",
   572 => x"2daee008",
   573 => x"aee00880",
   574 => x"fffffff8",
   575 => x"06555c73",
   576 => x"80ffffff",
   577 => x"f82e9238",
   578 => x"aee008fe",
   579 => x"05b38c08",
   580 => x"29b39c08",
   581 => x"055790b5",
   582 => x"04805473",
   583 => x"aee00c02",
   584 => x"b8050d04",
   585 => x"02f4050d",
   586 => x"74700881",
   587 => x"05710c70",
   588 => x"08b39008",
   589 => x"06535371",
   590 => x"8e388813",
   591 => x"08518f9e",
   592 => x"2daee008",
   593 => x"88140c81",
   594 => x"0baee00c",
   595 => x"028c050d",
   596 => x"0402f005",
   597 => x"0d758811",
   598 => x"08fe05b3",
   599 => x"8c0829b3",
   600 => x"9c081172",
   601 => x"08b39008",
   602 => x"06057955",
   603 => x"53545498",
   604 => x"d62daee0",
   605 => x"0853aee0",
   606 => x"08802e83",
   607 => x"38815372",
   608 => x"aee00c02",
   609 => x"90050d04",
   610 => x"b39408ae",
   611 => x"e00c0402",
   612 => x"f4050dd4",
   613 => x"5281ff72",
   614 => x"0c710853",
   615 => x"81ff720c",
   616 => x"72882b83",
   617 => x"fe800672",
   618 => x"087081ff",
   619 => x"06515253",
   620 => x"81ff720c",
   621 => x"72710788",
   622 => x"2b720870",
   623 => x"81ff0651",
   624 => x"525381ff",
   625 => x"720c7271",
   626 => x"07882b72",
   627 => x"087081ff",
   628 => x"067207ae",
   629 => x"e00c5253",
   630 => x"028c050d",
   631 => x"0402f405",
   632 => x"0d747671",
   633 => x"81ff06d4",
   634 => x"0c5353b3",
   635 => x"bc088538",
   636 => x"71892b52",
   637 => x"71982ad4",
   638 => x"0c71902a",
   639 => x"7081ff06",
   640 => x"d40c5171",
   641 => x"882a7081",
   642 => x"ff06d40c",
   643 => x"517181ff",
   644 => x"06d40c72",
   645 => x"902a7081",
   646 => x"ff06d40c",
   647 => x"51d40870",
   648 => x"81ff0651",
   649 => x"5182b8bf",
   650 => x"527081ff",
   651 => x"2e098106",
   652 => x"943881ff",
   653 => x"0bd40cd4",
   654 => x"087081ff",
   655 => x"06ff1454",
   656 => x"515171e5",
   657 => x"3870aee0",
   658 => x"0c028c05",
   659 => x"0d0402fc",
   660 => x"050d81c7",
   661 => x"5181ff0b",
   662 => x"d40cff11",
   663 => x"51708025",
   664 => x"f4380284",
   665 => x"050d0402",
   666 => x"f0050d94",
   667 => x"ce2d819c",
   668 => x"9f538052",
   669 => x"87fc80f7",
   670 => x"5193dd2d",
   671 => x"aee00854",
   672 => x"aee00881",
   673 => x"2e098106",
   674 => x"a33881ff",
   675 => x"0bd40c82",
   676 => x"0a52849c",
   677 => x"80e95193",
   678 => x"dd2daee0",
   679 => x"088b3881",
   680 => x"ff0bd40c",
   681 => x"735395b2",
   682 => x"0494ce2d",
   683 => x"ff135372",
   684 => x"c13872ae",
   685 => x"e00c0290",
   686 => x"050d0402",
   687 => x"f4050d81",
   688 => x"ff0bd40c",
   689 => x"93538052",
   690 => x"87fc80c1",
   691 => x"5193dd2d",
   692 => x"aee0088b",
   693 => x"3881ff0b",
   694 => x"d40c8153",
   695 => x"95e80494",
   696 => x"ce2dff13",
   697 => x"5372df38",
   698 => x"72aee00c",
   699 => x"028c050d",
   700 => x"0402f005",
   701 => x"0d94ce2d",
   702 => x"83aa5284",
   703 => x"9c80c851",
   704 => x"93dd2dae",
   705 => x"e008812e",
   706 => x"09810692",
   707 => x"38938f2d",
   708 => x"aee00883",
   709 => x"ffff0653",
   710 => x"7283aa2e",
   711 => x"973895bb",
   712 => x"2d96af04",
   713 => x"815497b4",
   714 => x"04abc851",
   715 => x"85f02d80",
   716 => x"5497b404",
   717 => x"81ff0bd4",
   718 => x"0cb15394",
   719 => x"e72daee0",
   720 => x"08802e80",
   721 => x"e0388052",
   722 => x"87fc80fa",
   723 => x"5193dd2d",
   724 => x"aee00880",
   725 => x"c638aee0",
   726 => x"0852abe4",
   727 => x"519bf32d",
   728 => x"81ff0bd4",
   729 => x"0cd40870",
   730 => x"81ff0670",
   731 => x"54abf053",
   732 => x"51539bf3",
   733 => x"2d81ff0b",
   734 => x"d40c81ff",
   735 => x"0bd40c81",
   736 => x"ff0bd40c",
   737 => x"81ff0bd4",
   738 => x"0c72862a",
   739 => x"70810670",
   740 => x"56515372",
   741 => x"802e9d38",
   742 => x"96a404ae",
   743 => x"e00852ab",
   744 => x"e4519bf3",
   745 => x"2d72822e",
   746 => x"feff38ff",
   747 => x"135372ff",
   748 => x"8a387254",
   749 => x"73aee00c",
   750 => x"0290050d",
   751 => x"0402f405",
   752 => x"0d810bb3",
   753 => x"bc0cd008",
   754 => x"708f2a70",
   755 => x"81065151",
   756 => x"5372f338",
   757 => x"72d00c94",
   758 => x"ce2dd008",
   759 => x"708f2a70",
   760 => x"81065151",
   761 => x"5372f338",
   762 => x"810bd00c",
   763 => x"87538052",
   764 => x"84d480c0",
   765 => x"5193dd2d",
   766 => x"aee00881",
   767 => x"2e9a3872",
   768 => x"822e0981",
   769 => x"068c38ac",
   770 => x"805185f0",
   771 => x"2d805398",
   772 => x"cd04ff13",
   773 => x"5372d738",
   774 => x"95f12dae",
   775 => x"e008b3bc",
   776 => x"0caee008",
   777 => x"8b388152",
   778 => x"87fc80d0",
   779 => x"5193dd2d",
   780 => x"81ff0bd4",
   781 => x"0cd00870",
   782 => x"8f2a7081",
   783 => x"06515153",
   784 => x"72f33872",
   785 => x"d00c81ff",
   786 => x"0bd40c81",
   787 => x"5372aee0",
   788 => x"0c028c05",
   789 => x"0d0402e0",
   790 => x"050d797b",
   791 => x"57578058",
   792 => x"81ff0bd4",
   793 => x"0cd00870",
   794 => x"8f2a7081",
   795 => x"06515154",
   796 => x"73f33882",
   797 => x"810bd00c",
   798 => x"81ff0bd4",
   799 => x"0c765287",
   800 => x"fc80d151",
   801 => x"93dd2d80",
   802 => x"dbc6df55",
   803 => x"aee00880",
   804 => x"2e9038ae",
   805 => x"e0085376",
   806 => x"52ac9851",
   807 => x"9bf32d99",
   808 => x"f00481ff",
   809 => x"0bd40cd4",
   810 => x"087081ff",
   811 => x"06515473",
   812 => x"81fe2e09",
   813 => x"81069d38",
   814 => x"80ff5493",
   815 => x"8f2daee0",
   816 => x"08767084",
   817 => x"05580cff",
   818 => x"14547380",
   819 => x"25ed3881",
   820 => x"5899da04",
   821 => x"ff155574",
   822 => x"c93881ff",
   823 => x"0bd40cd0",
   824 => x"08708f2a",
   825 => x"70810651",
   826 => x"515473f3",
   827 => x"3873d00c",
   828 => x"77aee00c",
   829 => x"02a0050d",
   830 => x"04b3bc08",
   831 => x"aee00c04",
   832 => x"02e8050d",
   833 => x"80785755",
   834 => x"75708405",
   835 => x"57085380",
   836 => x"5472982a",
   837 => x"73882b54",
   838 => x"5271802e",
   839 => x"a238c008",
   840 => x"70882a70",
   841 => x"81065151",
   842 => x"5170802e",
   843 => x"f13871c0",
   844 => x"0c811581",
   845 => x"15555583",
   846 => x"7425d638",
   847 => x"71ca3874",
   848 => x"aee00c02",
   849 => x"98050d04",
   850 => x"02f4050d",
   851 => x"7470882a",
   852 => x"83fe8006",
   853 => x"7072982a",
   854 => x"0772882b",
   855 => x"87fc8080",
   856 => x"0673982b",
   857 => x"81f00a06",
   858 => x"71730707",
   859 => x"aee00c56",
   860 => x"51535102",
   861 => x"8c050d04",
   862 => x"02f8050d",
   863 => x"028e0580",
   864 => x"f52d7488",
   865 => x"2b077083",
   866 => x"ffff06ae",
   867 => x"e00c5102",
   868 => x"88050d04",
   869 => x"02ec050d",
   870 => x"76538055",
   871 => x"7275258b",
   872 => x"38ad5182",
   873 => x"ee2d7209",
   874 => x"81055372",
   875 => x"802eb538",
   876 => x"8754729c",
   877 => x"2a73842b",
   878 => x"54527180",
   879 => x"2e833881",
   880 => x"55897225",
   881 => x"8738b712",
   882 => x"529bcf04",
   883 => x"b0125274",
   884 => x"802e8638",
   885 => x"715182ee",
   886 => x"2dff1454",
   887 => x"738025d2",
   888 => x"389be904",
   889 => x"b05182ee",
   890 => x"2d800bae",
   891 => x"e00c0294",
   892 => x"050d0402",
   893 => x"c0050d02",
   894 => x"80c40557",
   895 => x"80707870",
   896 => x"84055a08",
   897 => x"72415f5d",
   898 => x"587c7084",
   899 => x"055e085a",
   900 => x"805b7998",
   901 => x"2a7a882b",
   902 => x"5b567586",
   903 => x"38775f9d",
   904 => x"eb047d80",
   905 => x"2e81a238",
   906 => x"805e7580",
   907 => x"e42e8a38",
   908 => x"7580f82e",
   909 => x"09810689",
   910 => x"38768418",
   911 => x"71085e58",
   912 => x"547580e4",
   913 => x"2e9f3875",
   914 => x"80e4268a",
   915 => x"387580e3",
   916 => x"2ebe389d",
   917 => x"9b047580",
   918 => x"f32ea338",
   919 => x"7580f82e",
   920 => x"89389d9b",
   921 => x"048a539c",
   922 => x"ec049053",
   923 => x"b3c0527b",
   924 => x"519b942d",
   925 => x"aee008b3",
   926 => x"c05a559d",
   927 => x"ab047684",
   928 => x"18710870",
   929 => x"545b5854",
   930 => x"9a802d80",
   931 => x"559dab04",
   932 => x"76841871",
   933 => x"08585854",
   934 => x"9dd604a5",
   935 => x"5182ee2d",
   936 => x"755182ee",
   937 => x"2d821858",
   938 => x"9dde0474",
   939 => x"ff165654",
   940 => x"807425aa",
   941 => x"38787081",
   942 => x"055a80f5",
   943 => x"2d705256",
   944 => x"82ee2d81",
   945 => x"18589dab",
   946 => x"0475a52e",
   947 => x"09810686",
   948 => x"38815e9d",
   949 => x"de047551",
   950 => x"82ee2d81",
   951 => x"1858811b",
   952 => x"5b837b25",
   953 => x"feac3875",
   954 => x"fe9f387e",
   955 => x"aee00c02",
   956 => x"80c0050d",
   957 => x"0402fc05",
   958 => x"0d725180",
   959 => x"710c800b",
   960 => x"84120c02",
   961 => x"84050d04",
   962 => x"02f0050d",
   963 => x"75700884",
   964 => x"12085353",
   965 => x"53ff5471",
   966 => x"712e9b38",
   967 => x"84130870",
   968 => x"8429148b",
   969 => x"1180f52d",
   970 => x"84160881",
   971 => x"11870684",
   972 => x"180c5256",
   973 => x"515173ae",
   974 => x"e00c0290",
   975 => x"050d0402",
   976 => x"f8050da1",
   977 => x"b62de008",
   978 => x"708b2a70",
   979 => x"81065152",
   980 => x"5270802e",
   981 => x"9d38b480",
   982 => x"08708429",
   983 => x"b4880573",
   984 => x"81ff0671",
   985 => x"0c5151b4",
   986 => x"80088111",
   987 => x"8706b480",
   988 => x"0c51800b",
   989 => x"b4a80ca1",
   990 => x"a92da1b0",
   991 => x"2d028805",
   992 => x"0d0402fc",
   993 => x"050da1b6",
   994 => x"2d810bb4",
   995 => x"a80ca1b0",
   996 => x"2db4a808",
   997 => x"5170fa38",
   998 => x"0284050d",
   999 => x"0402fc05",
  1000 => x"0db48051",
  1001 => x"9df52d9e",
  1002 => x"bf51a1a5",
  1003 => x"2da0cf2d",
  1004 => x"0284050d",
  1005 => x"0402f405",
  1006 => x"0da0b704",
  1007 => x"aee00881",
  1008 => x"f02e0981",
  1009 => x"06893881",
  1010 => x"0baed40c",
  1011 => x"a0b704ae",
  1012 => x"e00881e0",
  1013 => x"2e098106",
  1014 => x"8938810b",
  1015 => x"aed80ca0",
  1016 => x"b704aee0",
  1017 => x"0852aed8",
  1018 => x"08802e88",
  1019 => x"38aee008",
  1020 => x"81800552",
  1021 => x"71842c72",
  1022 => x"8f065353",
  1023 => x"aed40880",
  1024 => x"2e993872",
  1025 => x"8429ae94",
  1026 => x"05721381",
  1027 => x"712b7009",
  1028 => x"73080673",
  1029 => x"0c515353",
  1030 => x"a0ad0472",
  1031 => x"8429ae94",
  1032 => x"05721383",
  1033 => x"712b7208",
  1034 => x"07720c53",
  1035 => x"53800bae",
  1036 => x"d80c800b",
  1037 => x"aed40cb4",
  1038 => x"80519e88",
  1039 => x"2daee008",
  1040 => x"ff24fef8",
  1041 => x"38800bae",
  1042 => x"e00c028c",
  1043 => x"050d0402",
  1044 => x"f8050dae",
  1045 => x"94528f51",
  1046 => x"80727084",
  1047 => x"05540cff",
  1048 => x"11517080",
  1049 => x"25f23802",
  1050 => x"88050d04",
  1051 => x"02f0050d",
  1052 => x"7551a1b6",
  1053 => x"2d70822c",
  1054 => x"fc06ae94",
  1055 => x"1172109e",
  1056 => x"06710870",
  1057 => x"722a7083",
  1058 => x"0682742b",
  1059 => x"70097406",
  1060 => x"760c5451",
  1061 => x"56575351",
  1062 => x"53a1b02d",
  1063 => x"71aee00c",
  1064 => x"0290050d",
  1065 => x"0471980c",
  1066 => x"04ffb008",
  1067 => x"aee00c04",
  1068 => x"810bffb0",
  1069 => x"0c04800b",
  1070 => x"ffb00c04",
  1071 => x"02fc050d",
  1072 => x"800baedc",
  1073 => x"0c805184",
  1074 => x"e52d0284",
  1075 => x"050d0402",
  1076 => x"f0050db4",
  1077 => x"ac085481",
  1078 => x"f72d800b",
  1079 => x"b4b40c73",
  1080 => x"08802e80",
  1081 => x"eb38820b",
  1082 => x"aef40cb4",
  1083 => x"b4088f06",
  1084 => x"aef00c73",
  1085 => x"08527181",
  1086 => x"2ea43871",
  1087 => x"832e0981",
  1088 => x"06b93888",
  1089 => x"1480f52d",
  1090 => x"841508ac",
  1091 => x"b8535452",
  1092 => x"85f02d71",
  1093 => x"84291370",
  1094 => x"085252a2",
  1095 => x"bf04b4b0",
  1096 => x"08881508",
  1097 => x"2c708106",
  1098 => x"51527180",
  1099 => x"2e8738ac",
  1100 => x"bc51a2b8",
  1101 => x"04acc051",
  1102 => x"85f02d84",
  1103 => x"14085185",
  1104 => x"f02db4b4",
  1105 => x"088105b4",
  1106 => x"b40c8c14",
  1107 => x"54a1df04",
  1108 => x"0290050d",
  1109 => x"0471b4ac",
  1110 => x"0ca1cf2d",
  1111 => x"b4b408ff",
  1112 => x"05b4b80c",
  1113 => x"0402f005",
  1114 => x"0d8751a0",
  1115 => x"ec2daee0",
  1116 => x"08812a70",
  1117 => x"81065152",
  1118 => x"71802e8e",
  1119 => x"38aedc08",
  1120 => x"813270ae",
  1121 => x"dc0c5184",
  1122 => x"e52daedc",
  1123 => x"08802e82",
  1124 => x"9a3881f5",
  1125 => x"51a0ec2d",
  1126 => x"aee00881",
  1127 => x"2a708106",
  1128 => x"51527180",
  1129 => x"2e8f38b4",
  1130 => x"b8085271",
  1131 => x"802e8638",
  1132 => x"ff12b4b8",
  1133 => x"0c81f251",
  1134 => x"a0ec2dae",
  1135 => x"e008812a",
  1136 => x"70810651",
  1137 => x"5271802e",
  1138 => x"9538b4b4",
  1139 => x"08ff05b4",
  1140 => x"b8085452",
  1141 => x"72722586",
  1142 => x"388113b4",
  1143 => x"b80c80da",
  1144 => x"51a0ec2d",
  1145 => x"aee00881",
  1146 => x"2a708106",
  1147 => x"51527180",
  1148 => x"2e80fb38",
  1149 => x"b4ac08b4",
  1150 => x"b8085553",
  1151 => x"73802e8a",
  1152 => x"388c13ff",
  1153 => x"155553a3",
  1154 => x"fc047208",
  1155 => x"5271822e",
  1156 => x"a6387182",
  1157 => x"26893871",
  1158 => x"812ea538",
  1159 => x"a4ee0471",
  1160 => x"832ead38",
  1161 => x"71842e09",
  1162 => x"810680c2",
  1163 => x"38881308",
  1164 => x"51a2d52d",
  1165 => x"a4ee0488",
  1166 => x"13085271",
  1167 => x"2da4ee04",
  1168 => x"810b8814",
  1169 => x"082bb4b0",
  1170 => x"0832b4b0",
  1171 => x"0ca4eb04",
  1172 => x"881380f5",
  1173 => x"2d81058b",
  1174 => x"1480f52d",
  1175 => x"53547174",
  1176 => x"24833880",
  1177 => x"54738814",
  1178 => x"81b72da1",
  1179 => x"cf2d8054",
  1180 => x"800baef4",
  1181 => x"0c738f06",
  1182 => x"aef00ca0",
  1183 => x"5273b4b8",
  1184 => x"082e0981",
  1185 => x"069838b4",
  1186 => x"b408ff05",
  1187 => x"74327009",
  1188 => x"81057072",
  1189 => x"079f2a91",
  1190 => x"71315151",
  1191 => x"53537151",
  1192 => x"82ee2d81",
  1193 => x"14548e74",
  1194 => x"25c63802",
  1195 => x"90050d04",
  1196 => x"00ffffff",
  1197 => x"ff00ffff",
  1198 => x"ffff00ff",
  1199 => x"ffffff00",
  1200 => x"44495020",
  1201 => x"53776974",
  1202 => x"63686573",
  1203 => x"20100000",
  1204 => x"52657365",
  1205 => x"74000000",
  1206 => x"45786974",
  1207 => x"00000000",
  1208 => x"53442043",
  1209 => x"61726400",
  1210 => x"4a617061",
  1211 => x"6e657365",
  1212 => x"206b6579",
  1213 => x"626f6172",
  1214 => x"64206c61",
  1215 => x"796f7574",
  1216 => x"00000000",
  1217 => x"54757262",
  1218 => x"6f202831",
  1219 => x"302e3734",
  1220 => x"4d487a29",
  1221 => x"00000000",
  1222 => x"4261636b",
  1223 => x"00000000",
  1224 => x"32303438",
  1225 => x"4c422052",
  1226 => x"414d0000",
  1227 => x"34303936",
  1228 => x"4b422052",
  1229 => x"414d0000",
  1230 => x"536c323a",
  1231 => x"204e6f6e",
  1232 => x"65000000",
  1233 => x"536c323a",
  1234 => x"20455345",
  1235 => x"2d534343",
  1236 => x"20314d42",
  1237 => x"2f534343",
  1238 => x"2d490000",
  1239 => x"536c323a",
  1240 => x"20455345",
  1241 => x"2d52414d",
  1242 => x"20314d42",
  1243 => x"2f415343",
  1244 => x"49493800",
  1245 => x"536c323a",
  1246 => x"20455345",
  1247 => x"2d52414d",
  1248 => x"20314d42",
  1249 => x"2f415343",
  1250 => x"49493136",
  1251 => x"00000000",
  1252 => x"536c313a",
  1253 => x"204e6f6e",
  1254 => x"65000000",
  1255 => x"536c313a",
  1256 => x"20455345",
  1257 => x"2d534343",
  1258 => x"20314d42",
  1259 => x"2f534343",
  1260 => x"2d490000",
  1261 => x"536c313a",
  1262 => x"204d6567",
  1263 => x"6152414d",
  1264 => x"00000000",
  1265 => x"56474120",
  1266 => x"2d203331",
  1267 => x"4b487a2c",
  1268 => x"20363048",
  1269 => x"7a000000",
  1270 => x"56474120",
  1271 => x"2d203331",
  1272 => x"4b487a2c",
  1273 => x"20353048",
  1274 => x"7a000000",
  1275 => x"53434152",
  1276 => x"54202d20",
  1277 => x"31354b48",
  1278 => x"7a2c2035",
  1279 => x"30487a20",
  1280 => x"52474200",
  1281 => x"54562f53",
  1282 => x"6f756e64",
  1283 => x"202d2031",
  1284 => x"35487a00",
  1285 => x"496e6974",
  1286 => x"69616c69",
  1287 => x"7a696e67",
  1288 => x"20534420",
  1289 => x"63617264",
  1290 => x"0a000000",
  1291 => x"53444843",
  1292 => x"20636172",
  1293 => x"64206465",
  1294 => x"74656374",
  1295 => x"65642062",
  1296 => x"7574206e",
  1297 => x"6f740a73",
  1298 => x"7570706f",
  1299 => x"72746564",
  1300 => x"202d2064",
  1301 => x"69736162",
  1302 => x"6c696e67",
  1303 => x"20534420",
  1304 => x"63617264",
  1305 => x"0a10204f",
  1306 => x"4b0a0000",
  1307 => x"46617433",
  1308 => x"32206669",
  1309 => x"6c657379",
  1310 => x"7374656d",
  1311 => x"20646574",
  1312 => x"65637465",
  1313 => x"64206275",
  1314 => x"74206e6f",
  1315 => x"740a7375",
  1316 => x"70706f72",
  1317 => x"74656420",
  1318 => x"2d206469",
  1319 => x"7361626c",
  1320 => x"696e6720",
  1321 => x"53442063",
  1322 => x"6172640a",
  1323 => x"10204f4b",
  1324 => x"0a000000",
  1325 => x"54727969",
  1326 => x"6e67204d",
  1327 => x"53583342",
  1328 => x"494f532e",
  1329 => x"5359532e",
  1330 => x"2e2e0a00",
  1331 => x"4d535833",
  1332 => x"42494f53",
  1333 => x"53595300",
  1334 => x"54727969",
  1335 => x"6e672042",
  1336 => x"494f535f",
  1337 => x"4d32502e",
  1338 => x"524f4d2e",
  1339 => x"2e2e0a00",
  1340 => x"42494f53",
  1341 => x"5f4d3250",
  1342 => x"524f4d00",
  1343 => x"4f70656e",
  1344 => x"65642042",
  1345 => x"494f532c",
  1346 => x"206c6f61",
  1347 => x"64696e67",
  1348 => x"2e2e2e0a",
  1349 => x"00000000",
  1350 => x"52656164",
  1351 => x"20626c6f",
  1352 => x"636b2066",
  1353 => x"61696c65",
  1354 => x"640a0000",
  1355 => x"4c6f6164",
  1356 => x"696e6720",
  1357 => x"42494f53",
  1358 => x"20666169",
  1359 => x"6c65640a",
  1360 => x"00000000",
  1361 => x"52656164",
  1362 => x"206f6620",
  1363 => x"4d425220",
  1364 => x"6661696c",
  1365 => x"65640a00",
  1366 => x"46415431",
  1367 => x"36202020",
  1368 => x"00000000",
  1369 => x"46415433",
  1370 => x"32202020",
  1371 => x"00000000",
  1372 => x"25642070",
  1373 => x"61727469",
  1374 => x"74696f6e",
  1375 => x"7320666f",
  1376 => x"756e640a",
  1377 => x"00000000",
  1378 => x"4e6f2070",
  1379 => x"61727469",
  1380 => x"74696f6e",
  1381 => x"20736967",
  1382 => x"6e617475",
  1383 => x"72652066",
  1384 => x"6f756e64",
  1385 => x"0a000000",
  1386 => x"556e7375",
  1387 => x"70706f72",
  1388 => x"74656420",
  1389 => x"70617274",
  1390 => x"6974696f",
  1391 => x"6e207479",
  1392 => x"7065210a",
  1393 => x"00000000",
  1394 => x"53444843",
  1395 => x"20496e69",
  1396 => x"7469616c",
  1397 => x"697a6174",
  1398 => x"696f6e20",
  1399 => x"6572726f",
  1400 => x"72210a00",
  1401 => x"434d4435",
  1402 => x"38202564",
  1403 => x"0a202000",
  1404 => x"434d4435",
  1405 => x"385f3220",
  1406 => x"25640a20",
  1407 => x"20000000",
  1408 => x"53442063",
  1409 => x"61726420",
  1410 => x"72657365",
  1411 => x"74206661",
  1412 => x"696c6564",
  1413 => x"210a0000",
  1414 => x"52656164",
  1415 => x"20636f6d",
  1416 => x"6d616e64",
  1417 => x"20666169",
  1418 => x"6c656420",
  1419 => x"61742025",
  1420 => x"64202825",
  1421 => x"64290a00",
  1422 => x"16200000",
  1423 => x"14200000",
  1424 => x"15200000",
  1425 => x"00000004",
  1426 => x"000012c0",
  1427 => x"00001674",
  1428 => x"00000002",
  1429 => x"000012d0",
  1430 => x"00000311",
  1431 => x"00000002",
  1432 => x"000012d8",
  1433 => x"000010bc",
  1434 => x"00000000",
  1435 => x"00000000",
  1436 => x"00000000",
  1437 => x"00000003",
  1438 => x"00001704",
  1439 => x"00000004",
  1440 => x"00000001",
  1441 => x"000012e0",
  1442 => x"00000002",
  1443 => x"00000003",
  1444 => x"000016f8",
  1445 => x"00000003",
  1446 => x"00000003",
  1447 => x"000016e8",
  1448 => x"00000004",
  1449 => x"00000001",
  1450 => x"000012e8",
  1451 => x"00000006",
  1452 => x"00000001",
  1453 => x"00001304",
  1454 => x"00000007",
  1455 => x"00000003",
  1456 => x"000016e0",
  1457 => x"00000002",
  1458 => x"00000004",
  1459 => x"00001318",
  1460 => x"00001644",
  1461 => x"00000000",
  1462 => x"00000000",
  1463 => x"00000000",
  1464 => x"00001320",
  1465 => x"0000132c",
  1466 => x"00001338",
  1467 => x"00001344",
  1468 => x"0000135c",
  1469 => x"00001374",
  1470 => x"00001390",
  1471 => x"0000139c",
  1472 => x"000013b4",
  1473 => x"000013c4",
  1474 => x"000013d8",
  1475 => x"000013ec",
  1476 => x"00001404",
  1477 => x"00000000",
  1478 => x"00000000",
  1479 => x"00000000",
  1480 => x"00000000",
  1481 => x"00000000",
  1482 => x"00000000",
  1483 => x"00000000",
  1484 => x"00000000",
  1485 => x"00000000",
  1486 => x"00000000",
  1487 => x"00000000",
  1488 => x"00000000",
  1489 => x"00000000",
  1490 => x"00000000",
  1491 => x"00000000",
  1492 => x"00000000",
  1493 => x"00000000",
  1494 => x"00000000",
  1495 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

