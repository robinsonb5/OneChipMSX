-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b0bb2",
     9 => x"f8080b0b",
    10 => x"0bb2fc08",
    11 => x"0b0b0bb3",
    12 => x"80080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"b3800c0b",
    16 => x"0b0bb2fc",
    17 => x"0c0b0b0b",
    18 => x"b2f80c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0ba3a4",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"b2f870b9",
    57 => x"d4278b38",
    58 => x"80717084",
    59 => x"05530c81",
    60 => x"e2048c51",
    61 => x"81f70402",
    62 => x"d8050d81",
    63 => x"0bfec40c",
    64 => x"b90bfec0",
    65 => x"0c840bfe",
    66 => x"c40ca3b4",
    67 => x"5195d02d",
    68 => x"92f12db2",
    69 => x"f808802e",
    70 => x"81b338a3",
    71 => x"cc5195d0",
    72 => x"2d84b02d",
    73 => x"a3e452b4",
    74 => x"b0518b95",
    75 => x"2db2f808",
    76 => x"81ff0653",
    77 => x"72802e81",
    78 => x"8e38a3f0",
    79 => x"5195d02d",
    80 => x"b4b40883",
    81 => x"ff05892a",
    82 => x"59805877",
    83 => x"792580fd",
    84 => x"38b4c852",
    85 => x"b4b0518d",
    86 => x"f02db2f8",
    87 => x"0881ff06",
    88 => x"5372802e",
    89 => x"80ca38b4",
    90 => x"c85a7785",
    91 => x"3877fec8",
    92 => x"0c83fc57",
    93 => x"79708405",
    94 => x"5b087082",
    95 => x"80297131",
    96 => x"71882c70",
    97 => x"81ff0673",
    98 => x"902c7081",
    99 => x"ff067598",
   100 => x"2afec80c",
   101 => x"fec80c58",
   102 => x"fec80c57",
   103 => x"fec80c53",
   104 => x"ab5195ae",
   105 => x"2dfc1757",
   106 => x"768025c8",
   107 => x"3883b604",
   108 => x"a48c5195",
   109 => x"d02db4b0",
   110 => x"518dc32d",
   111 => x"811858ae",
   112 => x"5195ae2d",
   113 => x"82cb04a4",
   114 => x"a05195d0",
   115 => x"2d800bfe",
   116 => x"c40ca4b8",
   117 => x"5195d02d",
   118 => x"9ef92da2",
   119 => x"a72d9f91",
   120 => x"2db2f808",
   121 => x"802ef738",
   122 => x"b2f80851",
   123 => x"95ae2d83",
   124 => x"de0402e8",
   125 => x"050d7779",
   126 => x"7b585555",
   127 => x"80537276",
   128 => x"25a33874",
   129 => x"70810556",
   130 => x"80f52d74",
   131 => x"70810556",
   132 => x"80f52d52",
   133 => x"5271712e",
   134 => x"86388151",
   135 => x"84a70481",
   136 => x"135383fe",
   137 => x"04805170",
   138 => x"b2f80c02",
   139 => x"98050d04",
   140 => x"02d8050d",
   141 => x"ff0bb8d0",
   142 => x"0c800bb8",
   143 => x"e40ca4d8",
   144 => x"5195d02d",
   145 => x"b4c85280",
   146 => x"51948b2d",
   147 => x"b2f80854",
   148 => x"b2f8088c",
   149 => x"38a4e851",
   150 => x"95d02d73",
   151 => x"558a8804",
   152 => x"a4fc5195",
   153 => x"d02d8056",
   154 => x"810bb4bc",
   155 => x"0c8853a5",
   156 => x"9452b4fe",
   157 => x"5183f22d",
   158 => x"b2f80876",
   159 => x"2e098106",
   160 => x"8738b2f8",
   161 => x"08b4bc0c",
   162 => x"8853a5a0",
   163 => x"52b59a51",
   164 => x"83f22db2",
   165 => x"f8088738",
   166 => x"b2f808b4",
   167 => x"bc0cb4bc",
   168 => x"0852a5ac",
   169 => x"5197d82d",
   170 => x"b4bc0880",
   171 => x"2e818738",
   172 => x"b88e0b80",
   173 => x"f52db88f",
   174 => x"0b80f52d",
   175 => x"71982b71",
   176 => x"902b07b8",
   177 => x"900b80f5",
   178 => x"2d70882b",
   179 => x"7207b891",
   180 => x"0b80f52d",
   181 => x"7107b8c6",
   182 => x"0b80f52d",
   183 => x"b8c70b80",
   184 => x"f52d7188",
   185 => x"2b07535f",
   186 => x"54525a56",
   187 => x"57557381",
   188 => x"abaa2e09",
   189 => x"81068d38",
   190 => x"75519698",
   191 => x"2db2f808",
   192 => x"56869404",
   193 => x"7382d4d5",
   194 => x"2e8a38a5",
   195 => x"c05195d0",
   196 => x"2d87c904",
   197 => x"7552a5e0",
   198 => x"5197d82d",
   199 => x"b4c85275",
   200 => x"51948b2d",
   201 => x"b2f80855",
   202 => x"b2f80880",
   203 => x"2e83d938",
   204 => x"a5f85195",
   205 => x"d02da6a0",
   206 => x"5197d82d",
   207 => x"8853a5a0",
   208 => x"52b59a51",
   209 => x"83f22db2",
   210 => x"f8088938",
   211 => x"810bb8e4",
   212 => x"0c86ef04",
   213 => x"8853a594",
   214 => x"52b4fe51",
   215 => x"83f22db2",
   216 => x"f808802e",
   217 => x"8a38a6b8",
   218 => x"5197d82d",
   219 => x"87c904b8",
   220 => x"c60b80f5",
   221 => x"2d547380",
   222 => x"d52e0981",
   223 => x"0680ca38",
   224 => x"b8c70b80",
   225 => x"f52d5473",
   226 => x"81aa2e09",
   227 => x"8106ba38",
   228 => x"800bb4c8",
   229 => x"0b80f52d",
   230 => x"56547481",
   231 => x"e92e8338",
   232 => x"81547481",
   233 => x"eb2e8c38",
   234 => x"80557375",
   235 => x"2e098106",
   236 => x"82d638b4",
   237 => x"d30b80f5",
   238 => x"2d59788d",
   239 => x"38b4d40b",
   240 => x"80f52d54",
   241 => x"73822e86",
   242 => x"3880558a",
   243 => x"8804b4d5",
   244 => x"0b80f52d",
   245 => x"70b8ec0c",
   246 => x"ff1170b8",
   247 => x"e00c5452",
   248 => x"a6d85197",
   249 => x"d82db4d6",
   250 => x"0b80f52d",
   251 => x"b4d70b80",
   252 => x"f52d5676",
   253 => x"05758280",
   254 => x"290570b8",
   255 => x"d40cb4d8",
   256 => x"0b80f52d",
   257 => x"70b8cc0c",
   258 => x"b8e40859",
   259 => x"57587680",
   260 => x"2e81a538",
   261 => x"8853a5a0",
   262 => x"52b59a51",
   263 => x"83f22d78",
   264 => x"55b2f808",
   265 => x"81e238b8",
   266 => x"ec087084",
   267 => x"2bb8c80c",
   268 => x"70b8e80c",
   269 => x"b4ed0b80",
   270 => x"f52db4ec",
   271 => x"0b80f52d",
   272 => x"71828029",
   273 => x"05b4ee0b",
   274 => x"80f52d70",
   275 => x"84808029",
   276 => x"12b4ef0b",
   277 => x"80f52d70",
   278 => x"81800a29",
   279 => x"1270b4c0",
   280 => x"0cb8cc08",
   281 => x"7129b8d4",
   282 => x"080570b8",
   283 => x"f40cb4f5",
   284 => x"0b80f52d",
   285 => x"b4f40b80",
   286 => x"f52d7182",
   287 => x"802905b4",
   288 => x"f60b80f5",
   289 => x"2d708480",
   290 => x"802912b4",
   291 => x"f70b80f5",
   292 => x"2d70982b",
   293 => x"81f00a06",
   294 => x"720570b4",
   295 => x"c40cfe11",
   296 => x"7e297705",
   297 => x"b8dc0c52",
   298 => x"5752575d",
   299 => x"5751525f",
   300 => x"525c5757",
   301 => x"578a8604",
   302 => x"b4da0b80",
   303 => x"f52db4d9",
   304 => x"0b80f52d",
   305 => x"71828029",
   306 => x"0570b8c8",
   307 => x"0c70a029",
   308 => x"83ff0570",
   309 => x"892a70b8",
   310 => x"e80cb4df",
   311 => x"0b80f52d",
   312 => x"b4de0b80",
   313 => x"f52d7182",
   314 => x"80290570",
   315 => x"b4c00c7b",
   316 => x"71291e70",
   317 => x"b8dc0c7d",
   318 => x"b4c40c73",
   319 => x"05b8f40c",
   320 => x"555e5151",
   321 => x"55558155",
   322 => x"74b2f80c",
   323 => x"02a8050d",
   324 => x"0402ec05",
   325 => x"0d767087",
   326 => x"2c7180ff",
   327 => x"06575553",
   328 => x"b8e4088a",
   329 => x"3872882c",
   330 => x"7381ff06",
   331 => x"565473b8",
   332 => x"d0082ea6",
   333 => x"38b8d408",
   334 => x"1452a6fc",
   335 => x"5197d82d",
   336 => x"b4c852b8",
   337 => x"d4081451",
   338 => x"948b2db2",
   339 => x"f80853b2",
   340 => x"f808802e",
   341 => x"b73873b8",
   342 => x"d00cb8e4",
   343 => x"08802e98",
   344 => x"38748429",
   345 => x"b4c80570",
   346 => x"08525396",
   347 => x"982db2f8",
   348 => x"08f00a06",
   349 => x"558b8a04",
   350 => x"7410b4c8",
   351 => x"057080e0",
   352 => x"2d525396",
   353 => x"c82db2f8",
   354 => x"08557453",
   355 => x"72b2f80c",
   356 => x"0294050d",
   357 => x"0402c805",
   358 => x"0d7f615f",
   359 => x"5c8057ff",
   360 => x"0bb8d00c",
   361 => x"b4c408b8",
   362 => x"dc085758",
   363 => x"b8e40877",
   364 => x"2e8a38b8",
   365 => x"ec08842b",
   366 => x"598bc204",
   367 => x"b8e80884",
   368 => x"2b59805a",
   369 => x"79792781",
   370 => x"b638798f",
   371 => x"06a01858",
   372 => x"54739738",
   373 => x"7552a79c",
   374 => x"5197d82d",
   375 => x"b4c85275",
   376 => x"51811656",
   377 => x"948b2db4",
   378 => x"c8578077",
   379 => x"80f52d56",
   380 => x"5474742e",
   381 => x"83388154",
   382 => x"7481e52e",
   383 => x"80fb3881",
   384 => x"70750655",
   385 => x"5d73802e",
   386 => x"80ef388b",
   387 => x"1780f52d",
   388 => x"98065b7a",
   389 => x"80e33876",
   390 => x"5195d02d",
   391 => x"8b537d52",
   392 => x"765183f2",
   393 => x"2db2f808",
   394 => x"80cf389c",
   395 => x"17085196",
   396 => x"982db2f8",
   397 => x"08841d0c",
   398 => x"9a1780e0",
   399 => x"2d5196c8",
   400 => x"2db2f808",
   401 => x"b2f80888",
   402 => x"1e0cb2f8",
   403 => x"085555b8",
   404 => x"e408802e",
   405 => x"98389417",
   406 => x"80e02d51",
   407 => x"96c82db2",
   408 => x"f808902b",
   409 => x"83fff00a",
   410 => x"06701651",
   411 => x"5473881d",
   412 => x"0c7a7c0c",
   413 => x"7c548dba",
   414 => x"04811a5a",
   415 => x"8bc404b8",
   416 => x"e408802e",
   417 => x"b3387751",
   418 => x"8a912db2",
   419 => x"f808b2f8",
   420 => x"0853a7bc",
   421 => x"525897d8",
   422 => x"2d7780ff",
   423 => x"fffff806",
   424 => x"547380ff",
   425 => x"fffff82e",
   426 => x"8f38fe18",
   427 => x"b8ec0829",
   428 => x"b8f40805",
   429 => x"568bc204",
   430 => x"805473b2",
   431 => x"f80c02b8",
   432 => x"050d0402",
   433 => x"f4050d74",
   434 => x"70088105",
   435 => x"710c7008",
   436 => x"b8e00806",
   437 => x"5353718e",
   438 => x"38881308",
   439 => x"518a912d",
   440 => x"b2f80888",
   441 => x"140c810b",
   442 => x"b2f80c02",
   443 => x"8c050d04",
   444 => x"02f0050d",
   445 => x"75881108",
   446 => x"fe05b8ec",
   447 => x"0829b8f4",
   448 => x"08117208",
   449 => x"b8e00806",
   450 => x"05795553",
   451 => x"5454948b",
   452 => x"2db2f808",
   453 => x"53b2f808",
   454 => x"802e8338",
   455 => x"815372b2",
   456 => x"f80c0290",
   457 => x"050d0402",
   458 => x"f4050dd4",
   459 => x"5281ff72",
   460 => x"0c710853",
   461 => x"81ff720c",
   462 => x"72882b83",
   463 => x"fe800672",
   464 => x"087081ff",
   465 => x"06515253",
   466 => x"81ff720c",
   467 => x"72710788",
   468 => x"2b720870",
   469 => x"81ff0651",
   470 => x"525381ff",
   471 => x"720c7271",
   472 => x"07882b72",
   473 => x"087081ff",
   474 => x"067207b2",
   475 => x"f80c5253",
   476 => x"028c050d",
   477 => x"0402f405",
   478 => x"0d747671",
   479 => x"81ff06d4",
   480 => x"0c5353b8",
   481 => x"f8088538",
   482 => x"71892b52",
   483 => x"71982ad4",
   484 => x"0c71902a",
   485 => x"7081ff06",
   486 => x"d40c5171",
   487 => x"882a7081",
   488 => x"ff06d40c",
   489 => x"517181ff",
   490 => x"06d40c72",
   491 => x"902a7081",
   492 => x"ff06d40c",
   493 => x"51d40870",
   494 => x"81ff0651",
   495 => x"5182b8bf",
   496 => x"527081ff",
   497 => x"2e098106",
   498 => x"943881ff",
   499 => x"0bd40cd4",
   500 => x"087081ff",
   501 => x"06ff1454",
   502 => x"515171e5",
   503 => x"3870b2f8",
   504 => x"0c028c05",
   505 => x"0d0402fc",
   506 => x"050d81c7",
   507 => x"5181ff0b",
   508 => x"d40cff11",
   509 => x"51708025",
   510 => x"f4380284",
   511 => x"050d0402",
   512 => x"f0050d8f",
   513 => x"e62d819c",
   514 => x"9f538052",
   515 => x"87fc80f7",
   516 => x"518ef52d",
   517 => x"b2f80854",
   518 => x"b2f80881",
   519 => x"2e098106",
   520 => x"a33881ff",
   521 => x"0bd40c82",
   522 => x"0a52849c",
   523 => x"80e9518e",
   524 => x"f52db2f8",
   525 => x"088b3881",
   526 => x"ff0bd40c",
   527 => x"735390ca",
   528 => x"048fe62d",
   529 => x"ff135372",
   530 => x"c13872b2",
   531 => x"f80c0290",
   532 => x"050d0402",
   533 => x"f4050d81",
   534 => x"ff0bd40c",
   535 => x"a7d45195",
   536 => x"d02d9353",
   537 => x"805287fc",
   538 => x"80c1518e",
   539 => x"f52db2f8",
   540 => x"088b3881",
   541 => x"ff0bd40c",
   542 => x"81539186",
   543 => x"048fe62d",
   544 => x"ff135372",
   545 => x"df3872b2",
   546 => x"f80c028c",
   547 => x"050d0402",
   548 => x"f0050d8f",
   549 => x"e62d83aa",
   550 => x"52849c80",
   551 => x"c8518ef5",
   552 => x"2db2f808",
   553 => x"b2f80853",
   554 => x"a7e05253",
   555 => x"97d82d72",
   556 => x"812e0981",
   557 => x"069c388e",
   558 => x"a72db2f8",
   559 => x"0883ffff",
   560 => x"06537283",
   561 => x"aa2ea138",
   562 => x"b2f80852",
   563 => x"a7f85197",
   564 => x"d82d90d3",
   565 => x"2d91e304",
   566 => x"815492e8",
   567 => x"04a89051",
   568 => x"97d82d80",
   569 => x"5492e804",
   570 => x"81ff0bd4",
   571 => x"0cb1538f",
   572 => x"ff2db2f8",
   573 => x"08802e80",
   574 => x"e0388052",
   575 => x"87fc80fa",
   576 => x"518ef52d",
   577 => x"b2f80880",
   578 => x"c638b2f8",
   579 => x"0852a8ac",
   580 => x"5197d82d",
   581 => x"81ff0bd4",
   582 => x"0cd40870",
   583 => x"81ff0670",
   584 => x"54a8b853",
   585 => x"515397d8",
   586 => x"2d81ff0b",
   587 => x"d40c81ff",
   588 => x"0bd40c81",
   589 => x"ff0bd40c",
   590 => x"81ff0bd4",
   591 => x"0c72862a",
   592 => x"70810670",
   593 => x"56515372",
   594 => x"802e9d38",
   595 => x"91d804b2",
   596 => x"f80852a8",
   597 => x"ac5197d8",
   598 => x"2d72822e",
   599 => x"feff38ff",
   600 => x"135372ff",
   601 => x"8a387254",
   602 => x"73b2f80c",
   603 => x"0290050d",
   604 => x"0402f405",
   605 => x"0d810bb8",
   606 => x"f80cd008",
   607 => x"708f2a70",
   608 => x"81065151",
   609 => x"5372f338",
   610 => x"72d00c8f",
   611 => x"e62da8c8",
   612 => x"5195d02d",
   613 => x"d008708f",
   614 => x"2a708106",
   615 => x"51515372",
   616 => x"f338810b",
   617 => x"d00c8753",
   618 => x"805284d4",
   619 => x"80c0518e",
   620 => x"f52db2f8",
   621 => x"08812e94",
   622 => x"3872822e",
   623 => x"09810686",
   624 => x"38805393",
   625 => x"fc04ff13",
   626 => x"5372dd38",
   627 => x"918f2db2",
   628 => x"f808b8f8",
   629 => x"0c815287",
   630 => x"fc80d051",
   631 => x"8ef52d81",
   632 => x"ff0bd40c",
   633 => x"d008708f",
   634 => x"2a708106",
   635 => x"51515372",
   636 => x"f33872d0",
   637 => x"0c81ff0b",
   638 => x"d40c8153",
   639 => x"72b2f80c",
   640 => x"028c050d",
   641 => x"04800bb2",
   642 => x"f80c0402",
   643 => x"e0050d79",
   644 => x"7b575780",
   645 => x"5881ff0b",
   646 => x"d40cd008",
   647 => x"708f2a70",
   648 => x"81065151",
   649 => x"5473f338",
   650 => x"82810bd0",
   651 => x"0c81ff0b",
   652 => x"d40c7652",
   653 => x"87fc80d1",
   654 => x"518ef52d",
   655 => x"80dbc6df",
   656 => x"55b2f808",
   657 => x"802e9038",
   658 => x"b2f80853",
   659 => x"7652a8d4",
   660 => x"5197d82d",
   661 => x"95a50481",
   662 => x"ff0bd40c",
   663 => x"d4087081",
   664 => x"ff065154",
   665 => x"7381fe2e",
   666 => x"0981069d",
   667 => x"3880ff54",
   668 => x"8ea72db2",
   669 => x"f8087670",
   670 => x"8405580c",
   671 => x"ff145473",
   672 => x"8025ed38",
   673 => x"8158958f",
   674 => x"04ff1555",
   675 => x"74c93881",
   676 => x"ff0bd40c",
   677 => x"d008708f",
   678 => x"2a708106",
   679 => x"51515473",
   680 => x"f33873d0",
   681 => x"0c77b2f8",
   682 => x"0c02a005",
   683 => x"0d0402f8",
   684 => x"050d7352",
   685 => x"c0087088",
   686 => x"2a708106",
   687 => x"51515170",
   688 => x"802ef138",
   689 => x"71c00c71",
   690 => x"b2f80c02",
   691 => x"88050d04",
   692 => x"02e8050d",
   693 => x"80785755",
   694 => x"75708405",
   695 => x"57085380",
   696 => x"5472982a",
   697 => x"73882b54",
   698 => x"5271802e",
   699 => x"a238c008",
   700 => x"70882a70",
   701 => x"81065151",
   702 => x"5170802e",
   703 => x"f13871c0",
   704 => x"0c811581",
   705 => x"15555583",
   706 => x"7425d638",
   707 => x"71ca3874",
   708 => x"b2f80c02",
   709 => x"98050d04",
   710 => x"02f4050d",
   711 => x"7470882a",
   712 => x"83fe8006",
   713 => x"7072982a",
   714 => x"0772882b",
   715 => x"87fc8080",
   716 => x"0673982b",
   717 => x"81f00a06",
   718 => x"71730707",
   719 => x"b2f80c56",
   720 => x"51535102",
   721 => x"8c050d04",
   722 => x"02f8050d",
   723 => x"028e0580",
   724 => x"f52d7488",
   725 => x"2b077083",
   726 => x"ffff06b2",
   727 => x"f80c5102",
   728 => x"88050d04",
   729 => x"02f8050d",
   730 => x"7370902b",
   731 => x"71902a07",
   732 => x"b2f80c52",
   733 => x"0288050d",
   734 => x"0402ec05",
   735 => x"0d765380",
   736 => x"55727525",
   737 => x"8b38ad51",
   738 => x"95ae2d72",
   739 => x"09810553",
   740 => x"72802eb5",
   741 => x"38875472",
   742 => x"9c2a7384",
   743 => x"2b545271",
   744 => x"802e8338",
   745 => x"81558972",
   746 => x"258738b7",
   747 => x"125297b4",
   748 => x"04b01252",
   749 => x"74802e86",
   750 => x"38715195",
   751 => x"ae2dff14",
   752 => x"54738025",
   753 => x"d23897ce",
   754 => x"04b05195",
   755 => x"ae2d800b",
   756 => x"b2f80c02",
   757 => x"94050d04",
   758 => x"02c0050d",
   759 => x"0280c405",
   760 => x"57807078",
   761 => x"7084055a",
   762 => x"0872415f",
   763 => x"5d587c70",
   764 => x"84055e08",
   765 => x"5a805b79",
   766 => x"982a7a88",
   767 => x"2b5b5675",
   768 => x"8638775f",
   769 => x"99d0047d",
   770 => x"802e81a2",
   771 => x"38805e75",
   772 => x"80e42e8a",
   773 => x"387580f8",
   774 => x"2e098106",
   775 => x"89387684",
   776 => x"1871085e",
   777 => x"58547580",
   778 => x"e42e9f38",
   779 => x"7580e426",
   780 => x"8a387580",
   781 => x"e32ebe38",
   782 => x"99800475",
   783 => x"80f32ea3",
   784 => x"387580f8",
   785 => x"2e893899",
   786 => x"80048a53",
   787 => x"98d10490",
   788 => x"53b3d852",
   789 => x"7b5196f9",
   790 => x"2db2f808",
   791 => x"b3d85a55",
   792 => x"99900476",
   793 => x"84187108",
   794 => x"70545b58",
   795 => x"5495d02d",
   796 => x"80559990",
   797 => x"04768418",
   798 => x"71085858",
   799 => x"5499bb04",
   800 => x"a55195ae",
   801 => x"2d755195",
   802 => x"ae2d8218",
   803 => x"5899c304",
   804 => x"74ff1656",
   805 => x"54807425",
   806 => x"aa387870",
   807 => x"81055a80",
   808 => x"f52d7052",
   809 => x"5695ae2d",
   810 => x"81185899",
   811 => x"900475a5",
   812 => x"2e098106",
   813 => x"8638815e",
   814 => x"99c30475",
   815 => x"5195ae2d",
   816 => x"81185881",
   817 => x"1b5b837b",
   818 => x"25feac38",
   819 => x"75fe9f38",
   820 => x"7eb2f80c",
   821 => x"0280c005",
   822 => x"0d0402ec",
   823 => x"050d7655",
   824 => x"7480f52d",
   825 => x"5170802e",
   826 => x"81f238b4",
   827 => x"9c087082",
   828 => x"808029a8",
   829 => x"f40805b4",
   830 => x"98081151",
   831 => x"5252718f",
   832 => x"24de3874",
   833 => x"70810556",
   834 => x"80f52d52",
   835 => x"71802e81",
   836 => x"cb387188",
   837 => x"2e098106",
   838 => x"9c38800b",
   839 => x"b4980825",
   840 => x"b838ff11",
   841 => x"51a07181",
   842 => x"b72db498",
   843 => x"08ff05b4",
   844 => x"980c9b81",
   845 => x"04718a2e",
   846 => x"0981069d",
   847 => x"38b49c08",
   848 => x"8105b49c",
   849 => x"0c800bb4",
   850 => x"980cb49c",
   851 => x"08828080",
   852 => x"29a8f408",
   853 => x"05519b81",
   854 => x"04717170",
   855 => x"81055381",
   856 => x"b72db498",
   857 => x"088105b4",
   858 => x"980cb498",
   859 => x"08a02e09",
   860 => x"81068e38",
   861 => x"800bb498",
   862 => x"0cb49c08",
   863 => x"8105b49c",
   864 => x"0c8f0bb4",
   865 => x"9c082580",
   866 => x"c738a8f4",
   867 => x"08828080",
   868 => x"11715355",
   869 => x"5381ff52",
   870 => x"73708405",
   871 => x"55087170",
   872 => x"8405530c",
   873 => x"ff125271",
   874 => x"8025ed38",
   875 => x"88801351",
   876 => x"8f528071",
   877 => x"70840553",
   878 => x"0cff1252",
   879 => x"718025f2",
   880 => x"38800bb4",
   881 => x"980c8f0b",
   882 => x"b49c0c9e",
   883 => x"80801351",
   884 => x"8f0bb49c",
   885 => x"0825feab",
   886 => x"3899e004",
   887 => x"0294050d",
   888 => x"0402f405",
   889 => x"0d029305",
   890 => x"80f52d02",
   891 => x"8c0581b7",
   892 => x"2d800284",
   893 => x"05890581",
   894 => x"b72d028c",
   895 => x"05fc0551",
   896 => x"99da2d81",
   897 => x"0bb2f80c",
   898 => x"028c050d",
   899 => x"0402fc05",
   900 => x"0d725199",
   901 => x"da2d800b",
   902 => x"b2f80c02",
   903 => x"84050d04",
   904 => x"02f8050d",
   905 => x"a8f40852",
   906 => x"8ffc5180",
   907 => x"72708405",
   908 => x"540cfc11",
   909 => x"51708025",
   910 => x"f2380288",
   911 => x"050d0402",
   912 => x"fc050d72",
   913 => x"5180710c",
   914 => x"800b8412",
   915 => x"0c800b88",
   916 => x"120c800b",
   917 => x"8c120c02",
   918 => x"84050d04",
   919 => x"02f0050d",
   920 => x"75700884",
   921 => x"12085353",
   922 => x"53ff5471",
   923 => x"712e9b38",
   924 => x"84130870",
   925 => x"84291493",
   926 => x"1180f52d",
   927 => x"84160881",
   928 => x"11870684",
   929 => x"180c5256",
   930 => x"515173b2",
   931 => x"f80c0290",
   932 => x"050d0402",
   933 => x"f4050d74",
   934 => x"70088412",
   935 => x"08535353",
   936 => x"7072248f",
   937 => x"38720884",
   938 => x"14087171",
   939 => x"31525252",
   940 => x"9dc00472",
   941 => x"08841408",
   942 => x"71713188",
   943 => x"05525252",
   944 => x"71b2f80c",
   945 => x"028c050d",
   946 => x"0402f805",
   947 => x"0da2ad2d",
   948 => x"a2a02de0",
   949 => x"08708b2a",
   950 => x"70810651",
   951 => x"52527080",
   952 => x"2e9d38b9",
   953 => x"84087084",
   954 => x"29b99405",
   955 => x"7381ff06",
   956 => x"710c5151",
   957 => x"b9840881",
   958 => x"118706b9",
   959 => x"840c5171",
   960 => x"8a2a7081",
   961 => x"06515170",
   962 => x"802ea838",
   963 => x"b98c08b9",
   964 => x"90085252",
   965 => x"71712e9b",
   966 => x"38b98c08",
   967 => x"708429b9",
   968 => x"b4057008",
   969 => x"e00c5151",
   970 => x"b98c0881",
   971 => x"118706b9",
   972 => x"8c0c51a2",
   973 => x"a72d0288",
   974 => x"050d0402",
   975 => x"f4050d74",
   976 => x"538c1308",
   977 => x"81118706",
   978 => x"88150854",
   979 => x"51517171",
   980 => x"2eef38a2",
   981 => x"ad2d8c13",
   982 => x"08708429",
   983 => x"1477b012",
   984 => x"0c51518c",
   985 => x"13088111",
   986 => x"87068c15",
   987 => x"0c519dc9",
   988 => x"2da2a72d",
   989 => x"028c050d",
   990 => x"0402fc05",
   991 => x"0db98451",
   992 => x"9cbf2d9d",
   993 => x"c951a29c",
   994 => x"2da1d42d",
   995 => x"0284050d",
   996 => x"0402e405",
   997 => x"0d8057a1",
   998 => x"9f04b2f8",
   999 => x"0881f02e",
  1000 => x"09810689",
  1001 => x"38810bb4",
  1002 => x"a80ca19f",
  1003 => x"04b2f808",
  1004 => x"81e02e09",
  1005 => x"81068938",
  1006 => x"810bb4ac",
  1007 => x"0ca19f04",
  1008 => x"b2f80854",
  1009 => x"b4ac0880",
  1010 => x"2e8838b2",
  1011 => x"f8088180",
  1012 => x"0554b4a8",
  1013 => x"08819c38",
  1014 => x"830ba8f8",
  1015 => x"1581b72d",
  1016 => x"7480ff24",
  1017 => x"b138b4a4",
  1018 => x"08822a70",
  1019 => x"8106b4a0",
  1020 => x"0870872b",
  1021 => x"81800778",
  1022 => x"11822b51",
  1023 => x"56585154",
  1024 => x"738b3875",
  1025 => x"81802915",
  1026 => x"70822b51",
  1027 => x"53aaf813",
  1028 => x"08537281",
  1029 => x"b638800b",
  1030 => x"b4ac0c74",
  1031 => x"80d92e80",
  1032 => x"c7387480",
  1033 => x"d9248f38",
  1034 => x"74922ebc",
  1035 => x"387480d8",
  1036 => x"2e9338a1",
  1037 => x"9a047480",
  1038 => x"f72ea038",
  1039 => x"7480fe2e",
  1040 => x"8f38a19a",
  1041 => x"04b4a408",
  1042 => x"8432b4a4",
  1043 => x"0ca0e304",
  1044 => x"b4a40881",
  1045 => x"32b4a40c",
  1046 => x"a0e304b4",
  1047 => x"a4088232",
  1048 => x"b4a40c81",
  1049 => x"57a19a04",
  1050 => x"b4a00881",
  1051 => x"07b4a00c",
  1052 => x"a19a04a8",
  1053 => x"f81480f5",
  1054 => x"2d81fe06",
  1055 => x"5372a8f8",
  1056 => x"1581b72d",
  1057 => x"74922e8a",
  1058 => x"387480d9",
  1059 => x"2e098106",
  1060 => x"8938b4a0",
  1061 => x"08fe06b4",
  1062 => x"a00c800b",
  1063 => x"b4a80cb9",
  1064 => x"84519cdc",
  1065 => x"2db2f808",
  1066 => x"55b2f808",
  1067 => x"ff24fdea",
  1068 => x"3876802e",
  1069 => x"943881ed",
  1070 => x"52b98451",
  1071 => x"9ebb2db4",
  1072 => x"a40852b9",
  1073 => x"84519ebb",
  1074 => x"2d805372",
  1075 => x"b2f80c02",
  1076 => x"9c050d04",
  1077 => x"02fc050d",
  1078 => x"8051800b",
  1079 => x"a8f81281",
  1080 => x"b72d8111",
  1081 => x"5181ff71",
  1082 => x"25f03802",
  1083 => x"84050d04",
  1084 => x"02f4050d",
  1085 => x"7451a2ad",
  1086 => x"2da8f811",
  1087 => x"80f52d70",
  1088 => x"81ff0671",
  1089 => x"fd065254",
  1090 => x"5271a8f8",
  1091 => x"1281b72d",
  1092 => x"a2a72d72",
  1093 => x"b2f80c02",
  1094 => x"8c050d04",
  1095 => x"71980c04",
  1096 => x"ffb008b2",
  1097 => x"f80c0481",
  1098 => x"0bffb00c",
  1099 => x"04800bff",
  1100 => x"b00c04b3",
  1101 => x"840802b3",
  1102 => x"840cff3d",
  1103 => x"0d800bb3",
  1104 => x"8408fc05",
  1105 => x"0cb38408",
  1106 => x"88050881",
  1107 => x"06ff1170",
  1108 => x"0970b384",
  1109 => x"088c0508",
  1110 => x"06b38408",
  1111 => x"fc050811",
  1112 => x"b38408fc",
  1113 => x"050cb384",
  1114 => x"08880508",
  1115 => x"812ab384",
  1116 => x"0888050c",
  1117 => x"b384088c",
  1118 => x"050810b3",
  1119 => x"84088c05",
  1120 => x"0c515151",
  1121 => x"51b38408",
  1122 => x"88050880",
  1123 => x"2e8438ff",
  1124 => x"b439b384",
  1125 => x"08fc0508",
  1126 => x"70b2f80c",
  1127 => x"51833d0d",
  1128 => x"b3840c04",
  1129 => x"00ffffff",
  1130 => x"ff00ffff",
  1131 => x"ffff00ff",
  1132 => x"ffffff00",
  1133 => x"496e6974",
  1134 => x"69616c69",
  1135 => x"7a696e67",
  1136 => x"20534420",
  1137 => x"63617264",
  1138 => x"0a000000",
  1139 => x"48756e74",
  1140 => x"696e6720",
  1141 => x"666f7220",
  1142 => x"70617274",
  1143 => x"6974696f",
  1144 => x"6e0a0000",
  1145 => x"42494f53",
  1146 => x"5f4d3250",
  1147 => x"524f4d00",
  1148 => x"4f70656e",
  1149 => x"65642066",
  1150 => x"696c652c",
  1151 => x"206c6f61",
  1152 => x"64696e67",
  1153 => x"2e2e2e0a",
  1154 => x"00000000",
  1155 => x"52656164",
  1156 => x"20626c6f",
  1157 => x"636b2066",
  1158 => x"61696c65",
  1159 => x"640a0000",
  1160 => x"4c6f6164",
  1161 => x"696e6720",
  1162 => x"42494f53",
  1163 => x"20666169",
  1164 => x"6c65640a",
  1165 => x"00000000",
  1166 => x"496e6974",
  1167 => x"69616c69",
  1168 => x"73696e67",
  1169 => x"2050532f",
  1170 => x"3220696e",
  1171 => x"74657266",
  1172 => x"6163652e",
  1173 => x"2e2e0a00",
  1174 => x"52656164",
  1175 => x"696e6720",
  1176 => x"4d42520a",
  1177 => x"00000000",
  1178 => x"52656164",
  1179 => x"206f6620",
  1180 => x"4d425220",
  1181 => x"6661696c",
  1182 => x"65640a00",
  1183 => x"4d425220",
  1184 => x"73756363",
  1185 => x"65737366",
  1186 => x"756c6c79",
  1187 => x"20726561",
  1188 => x"640a0000",
  1189 => x"46415431",
  1190 => x"36202020",
  1191 => x"00000000",
  1192 => x"46415433",
  1193 => x"32202020",
  1194 => x"00000000",
  1195 => x"50617274",
  1196 => x"6974696f",
  1197 => x"6e636f75",
  1198 => x"6e742025",
  1199 => x"640a0000",
  1200 => x"4e6f2070",
  1201 => x"61727469",
  1202 => x"74696f6e",
  1203 => x"20736967",
  1204 => x"6e617475",
  1205 => x"72652066",
  1206 => x"6f756e64",
  1207 => x"0a000000",
  1208 => x"52656164",
  1209 => x"696e6720",
  1210 => x"626f6f74",
  1211 => x"20736563",
  1212 => x"746f7220",
  1213 => x"25640a00",
  1214 => x"52656164",
  1215 => x"20626f6f",
  1216 => x"74207365",
  1217 => x"63746f72",
  1218 => x"2066726f",
  1219 => x"6d206669",
  1220 => x"72737420",
  1221 => x"70617274",
  1222 => x"6974696f",
  1223 => x"6e0a0000",
  1224 => x"48756e74",
  1225 => x"696e6720",
  1226 => x"666f7220",
  1227 => x"66696c65",
  1228 => x"73797374",
  1229 => x"656d0a00",
  1230 => x"556e7375",
  1231 => x"70706f72",
  1232 => x"74656420",
  1233 => x"70617274",
  1234 => x"6974696f",
  1235 => x"6e207479",
  1236 => x"7065210d",
  1237 => x"00000000",
  1238 => x"436c7573",
  1239 => x"74657220",
  1240 => x"73697a65",
  1241 => x"3a202564",
  1242 => x"2c20436c",
  1243 => x"75737465",
  1244 => x"72206d61",
  1245 => x"736b2c20",
  1246 => x"25640a00",
  1247 => x"47657443",
  1248 => x"6c757374",
  1249 => x"65722072",
  1250 => x"65616469",
  1251 => x"6e672073",
  1252 => x"6563746f",
  1253 => x"72202564",
  1254 => x"0a000000",
  1255 => x"52656164",
  1256 => x"696e6720",
  1257 => x"64697265",
  1258 => x"63746f72",
  1259 => x"79207365",
  1260 => x"63746f72",
  1261 => x"2025640a",
  1262 => x"00000000",
  1263 => x"47657446",
  1264 => x"41544c69",
  1265 => x"6e6b2072",
  1266 => x"65747572",
  1267 => x"6e656420",
  1268 => x"25640a00",
  1269 => x"436d645f",
  1270 => x"696e6974",
  1271 => x"0a000000",
  1272 => x"636d645f",
  1273 => x"434d4438",
  1274 => x"20726573",
  1275 => x"706f6e73",
  1276 => x"653a2025",
  1277 => x"640a0000",
  1278 => x"434d4438",
  1279 => x"5f342072",
  1280 => x"6573706f",
  1281 => x"6e73653a",
  1282 => x"2025640a",
  1283 => x"00000000",
  1284 => x"53444843",
  1285 => x"20496e69",
  1286 => x"7469616c",
  1287 => x"697a6174",
  1288 => x"696f6e20",
  1289 => x"6572726f",
  1290 => x"72210a00",
  1291 => x"434d4435",
  1292 => x"38202564",
  1293 => x"0a202000",
  1294 => x"434d4435",
  1295 => x"385f3220",
  1296 => x"25640a20",
  1297 => x"20000000",
  1298 => x"53504920",
  1299 => x"496e6974",
  1300 => x"28290a00",
  1301 => x"52656164",
  1302 => x"20636f6d",
  1303 => x"6d616e64",
  1304 => x"20666169",
  1305 => x"6c656420",
  1306 => x"61742025",
  1307 => x"64202825",
  1308 => x"64290a00",
  1309 => x"ffffe000",
  1310 => x"00000000",
  1311 => x"00000000",
  1312 => x"00000000",
  1313 => x"00000000",
  1314 => x"00000000",
  1315 => x"00000000",
  1316 => x"00000000",
  1317 => x"00000000",
  1318 => x"00000000",
  1319 => x"00000000",
  1320 => x"00000000",
  1321 => x"00000000",
  1322 => x"00000000",
  1323 => x"00000000",
  1324 => x"00000000",
  1325 => x"00000000",
  1326 => x"00000000",
  1327 => x"00000000",
  1328 => x"00000000",
  1329 => x"00000000",
  1330 => x"00000000",
  1331 => x"00000000",
  1332 => x"00000000",
  1333 => x"00000000",
  1334 => x"00000000",
  1335 => x"00000000",
  1336 => x"00000000",
  1337 => x"00000000",
  1338 => x"00000000",
  1339 => x"00000000",
  1340 => x"00000000",
  1341 => x"00000000",
  1342 => x"00000000",
  1343 => x"00000000",
  1344 => x"00000000",
  1345 => x"00000000",
  1346 => x"00000000",
  1347 => x"00000000",
  1348 => x"00000000",
  1349 => x"00000000",
  1350 => x"00000000",
  1351 => x"00000000",
  1352 => x"00000000",
  1353 => x"00000000",
  1354 => x"00000000",
  1355 => x"00000000",
  1356 => x"00000000",
  1357 => x"00000000",
  1358 => x"00000000",
  1359 => x"00000000",
  1360 => x"00000000",
  1361 => x"00000000",
  1362 => x"00000000",
  1363 => x"00000000",
  1364 => x"00000000",
  1365 => x"00000000",
  1366 => x"00000000",
  1367 => x"00000000",
  1368 => x"00000000",
  1369 => x"00000000",
  1370 => x"00000000",
  1371 => x"00000000",
  1372 => x"00000000",
  1373 => x"00000000",
  1374 => x"00000000",
  1375 => x"00000000",
  1376 => x"00000000",
  1377 => x"00000000",
  1378 => x"00000000",
  1379 => x"00000000",
  1380 => x"00000000",
  1381 => x"00000000",
  1382 => x"00000000",
  1383 => x"00000000",
  1384 => x"00000000",
  1385 => x"00000000",
  1386 => x"00000000",
  1387 => x"00000009",
  1388 => x"00000000",
  1389 => x"00000000",
  1390 => x"00000000",
  1391 => x"00000000",
  1392 => x"00000000",
  1393 => x"00000000",
  1394 => x"00000000",
  1395 => x"00000071",
  1396 => x"00000031",
  1397 => x"00000000",
  1398 => x"00000000",
  1399 => x"00000000",
  1400 => x"0000007a",
  1401 => x"00000073",
  1402 => x"00000061",
  1403 => x"00000077",
  1404 => x"00000032",
  1405 => x"00000000",
  1406 => x"00000000",
  1407 => x"00000063",
  1408 => x"00000078",
  1409 => x"00000064",
  1410 => x"00000065",
  1411 => x"00000034",
  1412 => x"00000033",
  1413 => x"00000000",
  1414 => x"00000000",
  1415 => x"00000020",
  1416 => x"00000076",
  1417 => x"00000066",
  1418 => x"00000074",
  1419 => x"00000072",
  1420 => x"00000035",
  1421 => x"00000000",
  1422 => x"00000000",
  1423 => x"0000006e",
  1424 => x"00000062",
  1425 => x"00000068",
  1426 => x"00000067",
  1427 => x"00000079",
  1428 => x"00000036",
  1429 => x"00000000",
  1430 => x"00000000",
  1431 => x"00000000",
  1432 => x"0000006d",
  1433 => x"0000006a",
  1434 => x"00000075",
  1435 => x"00000037",
  1436 => x"00000038",
  1437 => x"00000000",
  1438 => x"00000000",
  1439 => x"0000002c",
  1440 => x"0000006b",
  1441 => x"00000069",
  1442 => x"0000006f",
  1443 => x"00000030",
  1444 => x"00000039",
  1445 => x"00000000",
  1446 => x"00000000",
  1447 => x"0000002e",
  1448 => x"0000002f",
  1449 => x"0000006c",
  1450 => x"0000003b",
  1451 => x"00000070",
  1452 => x"0000002d",
  1453 => x"00000000",
  1454 => x"00000000",
  1455 => x"00000000",
  1456 => x"00000027",
  1457 => x"00000000",
  1458 => x"0000005b",
  1459 => x"0000003d",
  1460 => x"00000000",
  1461 => x"00000000",
  1462 => x"00000000",
  1463 => x"00000000",
  1464 => x"0000000a",
  1465 => x"0000005d",
  1466 => x"00000000",
  1467 => x"00000023",
  1468 => x"00000000",
  1469 => x"00000000",
  1470 => x"00000000",
  1471 => x"00000000",
  1472 => x"00000000",
  1473 => x"00000000",
  1474 => x"00000000",
  1475 => x"00000000",
  1476 => x"00000008",
  1477 => x"00000000",
  1478 => x"00000000",
  1479 => x"00000031",
  1480 => x"00000000",
  1481 => x"00000034",
  1482 => x"00000037",
  1483 => x"00000000",
  1484 => x"00000000",
  1485 => x"00000000",
  1486 => x"00000030",
  1487 => x"0000002e",
  1488 => x"00000032",
  1489 => x"00000035",
  1490 => x"00000036",
  1491 => x"00000038",
  1492 => x"0000001b",
  1493 => x"00000000",
  1494 => x"00000000",
  1495 => x"0000002b",
  1496 => x"00000033",
  1497 => x"00000000",
  1498 => x"0000002a",
  1499 => x"00000039",
  1500 => x"00000000",
  1501 => x"00000000",
  1502 => x"00000000",
  1503 => x"00000000",
  1504 => x"00000000",
  1505 => x"00000000",
  1506 => x"00000000",
  1507 => x"00000000",
  1508 => x"00000000",
  1509 => x"00000000",
  1510 => x"00000000",
  1511 => x"00000000",
  1512 => x"00000000",
  1513 => x"00000000",
  1514 => x"00000000",
  1515 => x"00000008",
  1516 => x"00000000",
  1517 => x"00000000",
  1518 => x"00000000",
  1519 => x"00000000",
  1520 => x"00000000",
  1521 => x"00000000",
  1522 => x"00000000",
  1523 => x"00000051",
  1524 => x"00000021",
  1525 => x"00000000",
  1526 => x"00000000",
  1527 => x"00000000",
  1528 => x"0000005a",
  1529 => x"00000053",
  1530 => x"00000041",
  1531 => x"00000057",
  1532 => x"00000022",
  1533 => x"00000000",
  1534 => x"00000000",
  1535 => x"00000043",
  1536 => x"00000058",
  1537 => x"00000044",
  1538 => x"00000045",
  1539 => x"00000024",
  1540 => x"000000a3",
  1541 => x"00000000",
  1542 => x"00000000",
  1543 => x"00000020",
  1544 => x"00000056",
  1545 => x"00000046",
  1546 => x"00000054",
  1547 => x"00000052",
  1548 => x"00000025",
  1549 => x"00000000",
  1550 => x"00000000",
  1551 => x"0000004e",
  1552 => x"00000042",
  1553 => x"00000048",
  1554 => x"00000047",
  1555 => x"00000059",
  1556 => x"0000005e",
  1557 => x"00000000",
  1558 => x"00000000",
  1559 => x"00000000",
  1560 => x"0000004d",
  1561 => x"0000004a",
  1562 => x"00000055",
  1563 => x"00000026",
  1564 => x"0000002a",
  1565 => x"00000000",
  1566 => x"00000000",
  1567 => x"0000003c",
  1568 => x"0000004b",
  1569 => x"00000049",
  1570 => x"0000004f",
  1571 => x"00000029",
  1572 => x"00000028",
  1573 => x"00000000",
  1574 => x"00000000",
  1575 => x"0000003e",
  1576 => x"0000003f",
  1577 => x"0000004c",
  1578 => x"0000003a",
  1579 => x"00000050",
  1580 => x"0000005f",
  1581 => x"00000000",
  1582 => x"00000000",
  1583 => x"00000000",
  1584 => x"0000003f",
  1585 => x"00000000",
  1586 => x"0000007b",
  1587 => x"0000002b",
  1588 => x"00000000",
  1589 => x"00000000",
  1590 => x"00000000",
  1591 => x"00000000",
  1592 => x"0000000a",
  1593 => x"0000007d",
  1594 => x"00000000",
  1595 => x"0000007e",
  1596 => x"00000000",
  1597 => x"00000000",
  1598 => x"00000000",
  1599 => x"00000000",
  1600 => x"00000000",
  1601 => x"00000000",
  1602 => x"00000000",
  1603 => x"00000000",
  1604 => x"00000009",
  1605 => x"00000000",
  1606 => x"00000000",
  1607 => x"00000031",
  1608 => x"00000000",
  1609 => x"00000034",
  1610 => x"00000037",
  1611 => x"00000000",
  1612 => x"00000000",
  1613 => x"00000000",
  1614 => x"00000030",
  1615 => x"0000002e",
  1616 => x"00000032",
  1617 => x"00000035",
  1618 => x"00000036",
  1619 => x"00000038",
  1620 => x"0000001b",
  1621 => x"00000000",
  1622 => x"00000000",
  1623 => x"0000002b",
  1624 => x"00000033",
  1625 => x"00000000",
  1626 => x"0000002a",
  1627 => x"00000039",
  1628 => x"00000000",
  1629 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

