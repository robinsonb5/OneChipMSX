-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b0bb3",
     9 => x"fc080b0b",
    10 => x"0bb48008",
    11 => x"0b0b0bb4",
    12 => x"84080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"b4840c0b",
    16 => x"0b0bb480",
    17 => x"0c0b0b0b",
    18 => x"b3fc0c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0ba4a8",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"b3fc70ba",
    57 => x"d8278b38",
    58 => x"80717084",
    59 => x"05530c81",
    60 => x"e2048c51",
    61 => x"81f70402",
    62 => x"d8050d81",
    63 => x"0bfec40c",
    64 => x"b90bfec0",
    65 => x"0c840bfe",
    66 => x"c40ca4b8",
    67 => x"5195eb2d",
    68 => x"9f942da2",
    69 => x"c22da4d8",
    70 => x"5195eb2d",
    71 => x"938c2db3",
    72 => x"fc08802e",
    73 => x"81ce38a4",
    74 => x"f05195eb",
    75 => x"2d84cb2d",
    76 => x"a58852b5",
    77 => x"b4518bb0",
    78 => x"2db3fc08",
    79 => x"81ff0653",
    80 => x"72802e81",
    81 => x"a938a594",
    82 => x"5195eb2d",
    83 => x"b5b80857",
    84 => x"805a7977",
    85 => x"25819d38",
    86 => x"9fac2db3",
    87 => x"fc08802e",
    88 => x"f738b5cc",
    89 => x"52b5b451",
    90 => x"8e8b2db3",
    91 => x"fc0881ff",
    92 => x"06537280",
    93 => x"2e80db38",
    94 => x"b5cc7a89",
    95 => x"2b53a7fc",
    96 => x"525997f3",
    97 => x"2d848052",
    98 => x"7851a2ce",
    99 => x"2d805883",
   100 => x"bf047870",
   101 => x"84055a08",
   102 => x"7081ff06",
   103 => x"71882c70",
   104 => x"81ff0673",
   105 => x"902c7081",
   106 => x"ff067598",
   107 => x"2afec80c",
   108 => x"fec80c58",
   109 => x"fec80c57",
   110 => x"fec80c84",
   111 => x"19595376",
   112 => x"53848077",
   113 => x"25843884",
   114 => x"80537278",
   115 => x"24c43883",
   116 => x"d804a5b0",
   117 => x"5195eb2d",
   118 => x"b5b4518d",
   119 => x"de2dfc80",
   120 => x"17811b5b",
   121 => x"57768024",
   122 => x"feee3883",
   123 => x"f404a5c4",
   124 => x"5195eb2d",
   125 => x"820bfec4",
   126 => x"0c9fac2d",
   127 => x"b3fc0880",
   128 => x"2ef738b3",
   129 => x"fc085195",
   130 => x"c92d83f9",
   131 => x"0402e805",
   132 => x"0d77797b",
   133 => x"58555580",
   134 => x"53727625",
   135 => x"a3387470",
   136 => x"81055680",
   137 => x"f52d7470",
   138 => x"81055680",
   139 => x"f52d5252",
   140 => x"71712e86",
   141 => x"38815184",
   142 => x"c2048113",
   143 => x"53849904",
   144 => x"805170b3",
   145 => x"fc0c0298",
   146 => x"050d0402",
   147 => x"d8050dff",
   148 => x"0bb9d40c",
   149 => x"800bb9e8",
   150 => x"0ca5dc51",
   151 => x"95eb2db5",
   152 => x"cc528051",
   153 => x"94a62db3",
   154 => x"fc0854b3",
   155 => x"fc088c38",
   156 => x"a5ec5195",
   157 => x"eb2d7355",
   158 => x"8aa304a6",
   159 => x"805195eb",
   160 => x"2d805681",
   161 => x"0bb5c00c",
   162 => x"8853a698",
   163 => x"52b68251",
   164 => x"848d2db3",
   165 => x"fc08762e",
   166 => x"09810687",
   167 => x"38b3fc08",
   168 => x"b5c00c88",
   169 => x"53a6a452",
   170 => x"b69e5184",
   171 => x"8d2db3fc",
   172 => x"088738b3",
   173 => x"fc08b5c0",
   174 => x"0cb5c008",
   175 => x"52a6b051",
   176 => x"97f32db5",
   177 => x"c008802e",
   178 => x"818738b9",
   179 => x"920b80f5",
   180 => x"2db9930b",
   181 => x"80f52d71",
   182 => x"982b7190",
   183 => x"2b07b994",
   184 => x"0b80f52d",
   185 => x"70882b72",
   186 => x"07b9950b",
   187 => x"80f52d71",
   188 => x"07b9ca0b",
   189 => x"80f52db9",
   190 => x"cb0b80f5",
   191 => x"2d71882b",
   192 => x"07535f54",
   193 => x"525a5657",
   194 => x"557381ab",
   195 => x"aa2e0981",
   196 => x"068d3875",
   197 => x"5196b32d",
   198 => x"b3fc0856",
   199 => x"86af0473",
   200 => x"82d4d52e",
   201 => x"8a38a6c4",
   202 => x"5195eb2d",
   203 => x"87e40475",
   204 => x"52a6e451",
   205 => x"97f32db5",
   206 => x"cc527551",
   207 => x"94a62db3",
   208 => x"fc0855b3",
   209 => x"fc08802e",
   210 => x"83d938a6",
   211 => x"fc5195eb",
   212 => x"2da7a451",
   213 => x"97f32d88",
   214 => x"53a6a452",
   215 => x"b69e5184",
   216 => x"8d2db3fc",
   217 => x"08893881",
   218 => x"0bb9e80c",
   219 => x"878a0488",
   220 => x"53a69852",
   221 => x"b6825184",
   222 => x"8d2db3fc",
   223 => x"08802e8a",
   224 => x"38a7bc51",
   225 => x"97f32d87",
   226 => x"e404b9ca",
   227 => x"0b80f52d",
   228 => x"547380d5",
   229 => x"2e098106",
   230 => x"80ca38b9",
   231 => x"cb0b80f5",
   232 => x"2d547381",
   233 => x"aa2e0981",
   234 => x"06ba3880",
   235 => x"0bb5cc0b",
   236 => x"80f52d56",
   237 => x"547481e9",
   238 => x"2e833881",
   239 => x"547481eb",
   240 => x"2e8c3880",
   241 => x"5573752e",
   242 => x"09810682",
   243 => x"d638b5d7",
   244 => x"0b80f52d",
   245 => x"59788d38",
   246 => x"b5d80b80",
   247 => x"f52d5473",
   248 => x"822e8638",
   249 => x"80558aa3",
   250 => x"04b5d90b",
   251 => x"80f52d70",
   252 => x"b9f00cff",
   253 => x"1170b9e4",
   254 => x"0c5452a7",
   255 => x"dc5197f3",
   256 => x"2db5da0b",
   257 => x"80f52db5",
   258 => x"db0b80f5",
   259 => x"2d567605",
   260 => x"75828029",
   261 => x"0570b9d8",
   262 => x"0cb5dc0b",
   263 => x"80f52d70",
   264 => x"b9d00cb9",
   265 => x"e8085957",
   266 => x"5876802e",
   267 => x"81a53888",
   268 => x"53a6a452",
   269 => x"b69e5184",
   270 => x"8d2d7855",
   271 => x"b3fc0881",
   272 => x"e238b9f0",
   273 => x"0870842b",
   274 => x"b9cc0c70",
   275 => x"b9ec0cb5",
   276 => x"f10b80f5",
   277 => x"2db5f00b",
   278 => x"80f52d71",
   279 => x"82802905",
   280 => x"b5f20b80",
   281 => x"f52d7084",
   282 => x"80802912",
   283 => x"b5f30b80",
   284 => x"f52d7081",
   285 => x"800a2912",
   286 => x"70b5c40c",
   287 => x"b9d00871",
   288 => x"29b9d808",
   289 => x"0570b9f8",
   290 => x"0cb5f90b",
   291 => x"80f52db5",
   292 => x"f80b80f5",
   293 => x"2d718280",
   294 => x"2905b5fa",
   295 => x"0b80f52d",
   296 => x"70848080",
   297 => x"2912b5fb",
   298 => x"0b80f52d",
   299 => x"70982b81",
   300 => x"f00a0672",
   301 => x"0570b5c8",
   302 => x"0cfe117e",
   303 => x"297705b9",
   304 => x"e00c5257",
   305 => x"52575d57",
   306 => x"51525f52",
   307 => x"5c575757",
   308 => x"8aa104b5",
   309 => x"de0b80f5",
   310 => x"2db5dd0b",
   311 => x"80f52d71",
   312 => x"82802905",
   313 => x"70b9cc0c",
   314 => x"70a02983",
   315 => x"ff057089",
   316 => x"2a70b9ec",
   317 => x"0cb5e30b",
   318 => x"80f52db5",
   319 => x"e20b80f5",
   320 => x"2d718280",
   321 => x"290570b5",
   322 => x"c40c7b71",
   323 => x"291e70b9",
   324 => x"e00c7db5",
   325 => x"c80c7305",
   326 => x"b9f80c55",
   327 => x"5e515155",
   328 => x"55815574",
   329 => x"b3fc0c02",
   330 => x"a8050d04",
   331 => x"02ec050d",
   332 => x"7670872c",
   333 => x"7180ff06",
   334 => x"575553b9",
   335 => x"e8088a38",
   336 => x"72882c73",
   337 => x"81ff0656",
   338 => x"5473b9d4",
   339 => x"082ea638",
   340 => x"b9d80814",
   341 => x"52a88051",
   342 => x"97f32db5",
   343 => x"cc52b9d8",
   344 => x"08145194",
   345 => x"a62db3fc",
   346 => x"0853b3fc",
   347 => x"08802eb7",
   348 => x"3873b9d4",
   349 => x"0cb9e808",
   350 => x"802e9838",
   351 => x"748429b5",
   352 => x"cc057008",
   353 => x"525396b3",
   354 => x"2db3fc08",
   355 => x"f00a0655",
   356 => x"8ba50474",
   357 => x"10b5cc05",
   358 => x"7080e02d",
   359 => x"525396e3",
   360 => x"2db3fc08",
   361 => x"55745372",
   362 => x"b3fc0c02",
   363 => x"94050d04",
   364 => x"02c8050d",
   365 => x"7f615f5c",
   366 => x"8057ff0b",
   367 => x"b9d40cb5",
   368 => x"c808b9e0",
   369 => x"085758b9",
   370 => x"e808772e",
   371 => x"8a38b9f0",
   372 => x"08842b59",
   373 => x"8bdd04b9",
   374 => x"ec08842b",
   375 => x"59805a79",
   376 => x"792781b6",
   377 => x"38798f06",
   378 => x"a0185854",
   379 => x"73973875",
   380 => x"52a8a051",
   381 => x"97f32db5",
   382 => x"cc527551",
   383 => x"81165694",
   384 => x"a62db5cc",
   385 => x"57807780",
   386 => x"f52d5654",
   387 => x"74742e83",
   388 => x"38815474",
   389 => x"81e52e80",
   390 => x"fb388170",
   391 => x"7506555d",
   392 => x"73802e80",
   393 => x"ef388b17",
   394 => x"80f52d98",
   395 => x"065b7a80",
   396 => x"e3387651",
   397 => x"95eb2d8b",
   398 => x"537d5276",
   399 => x"51848d2d",
   400 => x"b3fc0880",
   401 => x"cf389c17",
   402 => x"085196b3",
   403 => x"2db3fc08",
   404 => x"841d0c9a",
   405 => x"1780e02d",
   406 => x"5196e32d",
   407 => x"b3fc08b3",
   408 => x"fc08881e",
   409 => x"0cb3fc08",
   410 => x"5555b9e8",
   411 => x"08802e98",
   412 => x"38941780",
   413 => x"e02d5196",
   414 => x"e32db3fc",
   415 => x"08902b83",
   416 => x"fff00a06",
   417 => x"70165154",
   418 => x"73881d0c",
   419 => x"7a7c0c7c",
   420 => x"548dd504",
   421 => x"811a5a8b",
   422 => x"df04b9e8",
   423 => x"08802eb3",
   424 => x"3877518a",
   425 => x"ac2db3fc",
   426 => x"08b3fc08",
   427 => x"53a8c052",
   428 => x"5897f32d",
   429 => x"7780ffff",
   430 => x"fff80654",
   431 => x"7380ffff",
   432 => x"fff82e8f",
   433 => x"38fe18b9",
   434 => x"f00829b9",
   435 => x"f8080556",
   436 => x"8bdd0480",
   437 => x"5473b3fc",
   438 => x"0c02b805",
   439 => x"0d0402f4",
   440 => x"050d7470",
   441 => x"08810571",
   442 => x"0c7008b9",
   443 => x"e4080653",
   444 => x"53718e38",
   445 => x"88130851",
   446 => x"8aac2db3",
   447 => x"fc088814",
   448 => x"0c810bb3",
   449 => x"fc0c028c",
   450 => x"050d0402",
   451 => x"f0050d75",
   452 => x"881108fe",
   453 => x"05b9f008",
   454 => x"29b9f808",
   455 => x"117208b9",
   456 => x"e4080605",
   457 => x"79555354",
   458 => x"5494a62d",
   459 => x"b3fc0853",
   460 => x"b3fc0880",
   461 => x"2e833881",
   462 => x"5372b3fc",
   463 => x"0c029005",
   464 => x"0d0402f4",
   465 => x"050dd452",
   466 => x"81ff720c",
   467 => x"71085381",
   468 => x"ff720c72",
   469 => x"882b83fe",
   470 => x"80067208",
   471 => x"7081ff06",
   472 => x"51525381",
   473 => x"ff720c72",
   474 => x"7107882b",
   475 => x"72087081",
   476 => x"ff065152",
   477 => x"5381ff72",
   478 => x"0c727107",
   479 => x"882b7208",
   480 => x"7081ff06",
   481 => x"7207b3fc",
   482 => x"0c525302",
   483 => x"8c050d04",
   484 => x"02f4050d",
   485 => x"74767181",
   486 => x"ff06d40c",
   487 => x"5353b9fc",
   488 => x"08853871",
   489 => x"892b5271",
   490 => x"982ad40c",
   491 => x"71902a70",
   492 => x"81ff06d4",
   493 => x"0c517188",
   494 => x"2a7081ff",
   495 => x"06d40c51",
   496 => x"7181ff06",
   497 => x"d40c7290",
   498 => x"2a7081ff",
   499 => x"06d40c51",
   500 => x"d4087081",
   501 => x"ff065151",
   502 => x"82b8bf52",
   503 => x"7081ff2e",
   504 => x"09810694",
   505 => x"3881ff0b",
   506 => x"d40cd408",
   507 => x"7081ff06",
   508 => x"ff145451",
   509 => x"5171e538",
   510 => x"70b3fc0c",
   511 => x"028c050d",
   512 => x"0402fc05",
   513 => x"0d81c751",
   514 => x"81ff0bd4",
   515 => x"0cff1151",
   516 => x"708025f4",
   517 => x"38028405",
   518 => x"0d0402f0",
   519 => x"050d9081",
   520 => x"2d819c9f",
   521 => x"53805287",
   522 => x"fc80f751",
   523 => x"8f902db3",
   524 => x"fc0854b3",
   525 => x"fc08812e",
   526 => x"098106a3",
   527 => x"3881ff0b",
   528 => x"d40c820a",
   529 => x"52849c80",
   530 => x"e9518f90",
   531 => x"2db3fc08",
   532 => x"8b3881ff",
   533 => x"0bd40c73",
   534 => x"5390e504",
   535 => x"90812dff",
   536 => x"135372c1",
   537 => x"3872b3fc",
   538 => x"0c029005",
   539 => x"0d0402f4",
   540 => x"050d81ff",
   541 => x"0bd40ca8",
   542 => x"d85195eb",
   543 => x"2d935380",
   544 => x"5287fc80",
   545 => x"c1518f90",
   546 => x"2db3fc08",
   547 => x"8b3881ff",
   548 => x"0bd40c81",
   549 => x"5391a104",
   550 => x"90812dff",
   551 => x"135372df",
   552 => x"3872b3fc",
   553 => x"0c028c05",
   554 => x"0d0402f0",
   555 => x"050d9081",
   556 => x"2d83aa52",
   557 => x"849c80c8",
   558 => x"518f902d",
   559 => x"b3fc08b3",
   560 => x"fc0853a8",
   561 => x"e4525397",
   562 => x"f32d7281",
   563 => x"2e098106",
   564 => x"9c388ec2",
   565 => x"2db3fc08",
   566 => x"83ffff06",
   567 => x"537283aa",
   568 => x"2ea138b3",
   569 => x"fc0852a8",
   570 => x"fc5197f3",
   571 => x"2d90ee2d",
   572 => x"91fe0481",
   573 => x"54938304",
   574 => x"a9945197",
   575 => x"f32d8054",
   576 => x"93830481",
   577 => x"ff0bd40c",
   578 => x"b153909a",
   579 => x"2db3fc08",
   580 => x"802e80e0",
   581 => x"38805287",
   582 => x"fc80fa51",
   583 => x"8f902db3",
   584 => x"fc0880c6",
   585 => x"38b3fc08",
   586 => x"52a9b051",
   587 => x"97f32d81",
   588 => x"ff0bd40c",
   589 => x"d4087081",
   590 => x"ff067054",
   591 => x"a9bc5351",
   592 => x"5397f32d",
   593 => x"81ff0bd4",
   594 => x"0c81ff0b",
   595 => x"d40c81ff",
   596 => x"0bd40c81",
   597 => x"ff0bd40c",
   598 => x"72862a70",
   599 => x"81067056",
   600 => x"51537280",
   601 => x"2e9d3891",
   602 => x"f304b3fc",
   603 => x"0852a9b0",
   604 => x"5197f32d",
   605 => x"72822efe",
   606 => x"ff38ff13",
   607 => x"5372ff8a",
   608 => x"38725473",
   609 => x"b3fc0c02",
   610 => x"90050d04",
   611 => x"02f4050d",
   612 => x"810bb9fc",
   613 => x"0cd00870",
   614 => x"8f2a7081",
   615 => x"06515153",
   616 => x"72f33872",
   617 => x"d00c9081",
   618 => x"2da9cc51",
   619 => x"95eb2dd0",
   620 => x"08708f2a",
   621 => x"70810651",
   622 => x"515372f3",
   623 => x"38810bd0",
   624 => x"0c875380",
   625 => x"5284d480",
   626 => x"c0518f90",
   627 => x"2db3fc08",
   628 => x"812e9438",
   629 => x"72822e09",
   630 => x"81068638",
   631 => x"80539497",
   632 => x"04ff1353",
   633 => x"72dd3891",
   634 => x"aa2db3fc",
   635 => x"08b9fc0c",
   636 => x"815287fc",
   637 => x"80d0518f",
   638 => x"902d81ff",
   639 => x"0bd40cd0",
   640 => x"08708f2a",
   641 => x"70810651",
   642 => x"515372f3",
   643 => x"3872d00c",
   644 => x"81ff0bd4",
   645 => x"0c815372",
   646 => x"b3fc0c02",
   647 => x"8c050d04",
   648 => x"800bb3fc",
   649 => x"0c0402e0",
   650 => x"050d797b",
   651 => x"57578058",
   652 => x"81ff0bd4",
   653 => x"0cd00870",
   654 => x"8f2a7081",
   655 => x"06515154",
   656 => x"73f33882",
   657 => x"810bd00c",
   658 => x"81ff0bd4",
   659 => x"0c765287",
   660 => x"fc80d151",
   661 => x"8f902d80",
   662 => x"dbc6df55",
   663 => x"b3fc0880",
   664 => x"2e9038b3",
   665 => x"fc085376",
   666 => x"52a9d851",
   667 => x"97f32d95",
   668 => x"c00481ff",
   669 => x"0bd40cd4",
   670 => x"087081ff",
   671 => x"06515473",
   672 => x"81fe2e09",
   673 => x"81069d38",
   674 => x"80ff548e",
   675 => x"c22db3fc",
   676 => x"08767084",
   677 => x"05580cff",
   678 => x"14547380",
   679 => x"25ed3881",
   680 => x"5895aa04",
   681 => x"ff155574",
   682 => x"c93881ff",
   683 => x"0bd40cd0",
   684 => x"08708f2a",
   685 => x"70810651",
   686 => x"515473f3",
   687 => x"3873d00c",
   688 => x"77b3fc0c",
   689 => x"02a0050d",
   690 => x"0402f805",
   691 => x"0d7352c0",
   692 => x"0870882a",
   693 => x"70810651",
   694 => x"51517080",
   695 => x"2ef13871",
   696 => x"c00c71b3",
   697 => x"fc0c0288",
   698 => x"050d0402",
   699 => x"e8050d80",
   700 => x"78575575",
   701 => x"70840557",
   702 => x"08538054",
   703 => x"72982a73",
   704 => x"882b5452",
   705 => x"71802ea2",
   706 => x"38c00870",
   707 => x"882a7081",
   708 => x"06515151",
   709 => x"70802ef1",
   710 => x"3871c00c",
   711 => x"81158115",
   712 => x"55558374",
   713 => x"25d63871",
   714 => x"ca3874b3",
   715 => x"fc0c0298",
   716 => x"050d0402",
   717 => x"f4050d74",
   718 => x"70882a83",
   719 => x"fe800670",
   720 => x"72982a07",
   721 => x"72882b87",
   722 => x"fc808006",
   723 => x"73982b81",
   724 => x"f00a0671",
   725 => x"730707b3",
   726 => x"fc0c5651",
   727 => x"5351028c",
   728 => x"050d0402",
   729 => x"f8050d02",
   730 => x"8e0580f5",
   731 => x"2d74882b",
   732 => x"077083ff",
   733 => x"ff06b3fc",
   734 => x"0c510288",
   735 => x"050d0402",
   736 => x"f8050d73",
   737 => x"70902b71",
   738 => x"902a07b3",
   739 => x"fc0c5202",
   740 => x"88050d04",
   741 => x"02ec050d",
   742 => x"76538055",
   743 => x"7275258b",
   744 => x"38ad5195",
   745 => x"c92d7209",
   746 => x"81055372",
   747 => x"802eb538",
   748 => x"8754729c",
   749 => x"2a73842b",
   750 => x"54527180",
   751 => x"2e833881",
   752 => x"55897225",
   753 => x"8738b712",
   754 => x"5297cf04",
   755 => x"b0125274",
   756 => x"802e8638",
   757 => x"715195c9",
   758 => x"2dff1454",
   759 => x"738025d2",
   760 => x"3897e904",
   761 => x"b05195c9",
   762 => x"2d800bb3",
   763 => x"fc0c0294",
   764 => x"050d0402",
   765 => x"c0050d02",
   766 => x"80c40557",
   767 => x"80707870",
   768 => x"84055a08",
   769 => x"72415f5d",
   770 => x"587c7084",
   771 => x"055e085a",
   772 => x"805b7998",
   773 => x"2a7a882b",
   774 => x"5b567586",
   775 => x"38775f99",
   776 => x"eb047d80",
   777 => x"2e81a238",
   778 => x"805e7580",
   779 => x"e42e8a38",
   780 => x"7580f82e",
   781 => x"09810689",
   782 => x"38768418",
   783 => x"71085e58",
   784 => x"547580e4",
   785 => x"2e9f3875",
   786 => x"80e4268a",
   787 => x"387580e3",
   788 => x"2ebe3899",
   789 => x"9b047580",
   790 => x"f32ea338",
   791 => x"7580f82e",
   792 => x"8938999b",
   793 => x"048a5398",
   794 => x"ec049053",
   795 => x"b4dc527b",
   796 => x"5197942d",
   797 => x"b3fc08b4",
   798 => x"dc5a5599",
   799 => x"ab047684",
   800 => x"18710870",
   801 => x"545b5854",
   802 => x"95eb2d80",
   803 => x"5599ab04",
   804 => x"76841871",
   805 => x"08585854",
   806 => x"99d604a5",
   807 => x"5195c92d",
   808 => x"755195c9",
   809 => x"2d821858",
   810 => x"99de0474",
   811 => x"ff165654",
   812 => x"807425aa",
   813 => x"38787081",
   814 => x"055a80f5",
   815 => x"2d705256",
   816 => x"95c92d81",
   817 => x"185899ab",
   818 => x"0475a52e",
   819 => x"09810686",
   820 => x"38815e99",
   821 => x"de047551",
   822 => x"95c92d81",
   823 => x"1858811b",
   824 => x"5b837b25",
   825 => x"feac3875",
   826 => x"fe9f387e",
   827 => x"b3fc0c02",
   828 => x"80c0050d",
   829 => x"0402ec05",
   830 => x"0d765574",
   831 => x"80f52d51",
   832 => x"70802e81",
   833 => x"f238b5a0",
   834 => x"08708280",
   835 => x"8029a9f8",
   836 => x"0805b59c",
   837 => x"08115152",
   838 => x"52718f24",
   839 => x"de387470",
   840 => x"81055680",
   841 => x"f52d5271",
   842 => x"802e81cb",
   843 => x"3871882e",
   844 => x"0981069c",
   845 => x"38800bb5",
   846 => x"9c0825b8",
   847 => x"38ff1151",
   848 => x"a07181b7",
   849 => x"2db59c08",
   850 => x"ff05b59c",
   851 => x"0c9b9c04",
   852 => x"718a2e09",
   853 => x"81069d38",
   854 => x"b5a00881",
   855 => x"05b5a00c",
   856 => x"800bb59c",
   857 => x"0cb5a008",
   858 => x"82808029",
   859 => x"a9f80805",
   860 => x"519b9c04",
   861 => x"71717081",
   862 => x"055381b7",
   863 => x"2db59c08",
   864 => x"8105b59c",
   865 => x"0cb59c08",
   866 => x"a02e0981",
   867 => x"068e3880",
   868 => x"0bb59c0c",
   869 => x"b5a00881",
   870 => x"05b5a00c",
   871 => x"8f0bb5a0",
   872 => x"082580c7",
   873 => x"38a9f808",
   874 => x"82808011",
   875 => x"71535553",
   876 => x"81ff5273",
   877 => x"70840555",
   878 => x"08717084",
   879 => x"05530cff",
   880 => x"12527180",
   881 => x"25ed3888",
   882 => x"8013518f",
   883 => x"52807170",
   884 => x"8405530c",
   885 => x"ff125271",
   886 => x"8025f238",
   887 => x"800bb59c",
   888 => x"0c8f0bb5",
   889 => x"a00c9e80",
   890 => x"8013518f",
   891 => x"0bb5a008",
   892 => x"25feab38",
   893 => x"99fb0402",
   894 => x"94050d04",
   895 => x"02f4050d",
   896 => x"02930580",
   897 => x"f52d028c",
   898 => x"0581b72d",
   899 => x"80028405",
   900 => x"890581b7",
   901 => x"2d028c05",
   902 => x"fc055199",
   903 => x"f52d810b",
   904 => x"b3fc0c02",
   905 => x"8c050d04",
   906 => x"02fc050d",
   907 => x"725199f5",
   908 => x"2d800bb3",
   909 => x"fc0c0284",
   910 => x"050d0402",
   911 => x"f8050da9",
   912 => x"f808528f",
   913 => x"fc518072",
   914 => x"70840554",
   915 => x"0cfc1151",
   916 => x"708025f2",
   917 => x"38028805",
   918 => x"0d0402fc",
   919 => x"050d7251",
   920 => x"80710c80",
   921 => x"0b84120c",
   922 => x"800b8812",
   923 => x"0c800b8c",
   924 => x"120c0284",
   925 => x"050d0402",
   926 => x"f0050d75",
   927 => x"70088412",
   928 => x"08535353",
   929 => x"ff547171",
   930 => x"2e9b3884",
   931 => x"13087084",
   932 => x"29149311",
   933 => x"80f52d84",
   934 => x"16088111",
   935 => x"87068418",
   936 => x"0c525651",
   937 => x"5173b3fc",
   938 => x"0c029005",
   939 => x"0d0402f4",
   940 => x"050d7470",
   941 => x"08841208",
   942 => x"53535370",
   943 => x"72248f38",
   944 => x"72088414",
   945 => x"08717131",
   946 => x"5252529d",
   947 => x"db047208",
   948 => x"84140871",
   949 => x"71318805",
   950 => x"52525271",
   951 => x"b3fc0c02",
   952 => x"8c050d04",
   953 => x"02f8050d",
   954 => x"a2c82da2",
   955 => x"bb2de008",
   956 => x"708b2a70",
   957 => x"81065152",
   958 => x"5270802e",
   959 => x"9d38ba88",
   960 => x"08708429",
   961 => x"ba980573",
   962 => x"81ff0671",
   963 => x"0c5151ba",
   964 => x"88088111",
   965 => x"8706ba88",
   966 => x"0c51718a",
   967 => x"2a708106",
   968 => x"51517080",
   969 => x"2ea838ba",
   970 => x"9008ba94",
   971 => x"08525271",
   972 => x"712e9b38",
   973 => x"ba900870",
   974 => x"8429bab8",
   975 => x"057008e0",
   976 => x"0c5151ba",
   977 => x"90088111",
   978 => x"8706ba90",
   979 => x"0c51a2c2",
   980 => x"2d028805",
   981 => x"0d0402f4",
   982 => x"050d7453",
   983 => x"8c130881",
   984 => x"11870688",
   985 => x"15085451",
   986 => x"5171712e",
   987 => x"ef38a2c8",
   988 => x"2d8c1308",
   989 => x"70842914",
   990 => x"77b0120c",
   991 => x"51518c13",
   992 => x"08811187",
   993 => x"068c150c",
   994 => x"519de42d",
   995 => x"a2c22d02",
   996 => x"8c050d04",
   997 => x"02fc050d",
   998 => x"ba88519c",
   999 => x"da2d9de4",
  1000 => x"51a2b72d",
  1001 => x"a1ef2d02",
  1002 => x"84050d04",
  1003 => x"02e4050d",
  1004 => x"8057a1ba",
  1005 => x"04b3fc08",
  1006 => x"81f02e09",
  1007 => x"81068938",
  1008 => x"810bb5ac",
  1009 => x"0ca1ba04",
  1010 => x"b3fc0881",
  1011 => x"e02e0981",
  1012 => x"06893881",
  1013 => x"0bb5b00c",
  1014 => x"a1ba04b3",
  1015 => x"fc0854b5",
  1016 => x"b008802e",
  1017 => x"8838b3fc",
  1018 => x"08818005",
  1019 => x"54b5ac08",
  1020 => x"819c3883",
  1021 => x"0ba9fc15",
  1022 => x"81b72d74",
  1023 => x"80ff24b1",
  1024 => x"38b5a808",
  1025 => x"822a7081",
  1026 => x"06b5a408",
  1027 => x"70872b81",
  1028 => x"80077811",
  1029 => x"822b5156",
  1030 => x"58515473",
  1031 => x"8b387581",
  1032 => x"80291570",
  1033 => x"822b5153",
  1034 => x"abfc1308",
  1035 => x"537281b6",
  1036 => x"38800bb5",
  1037 => x"b00c7480",
  1038 => x"d92e80c7",
  1039 => x"387480d9",
  1040 => x"248f3874",
  1041 => x"922ebc38",
  1042 => x"7480d82e",
  1043 => x"9338a1b5",
  1044 => x"047480f7",
  1045 => x"2ea03874",
  1046 => x"80fe2e8f",
  1047 => x"38a1b504",
  1048 => x"b5a80884",
  1049 => x"32b5a80c",
  1050 => x"a0fe04b5",
  1051 => x"a8088132",
  1052 => x"b5a80ca0",
  1053 => x"fe04b5a8",
  1054 => x"088232b5",
  1055 => x"a80c8157",
  1056 => x"a1b504b5",
  1057 => x"a4088107",
  1058 => x"b5a40ca1",
  1059 => x"b504a9fc",
  1060 => x"1480f52d",
  1061 => x"81fe0653",
  1062 => x"72a9fc15",
  1063 => x"81b72d74",
  1064 => x"922e8a38",
  1065 => x"7480d92e",
  1066 => x"09810689",
  1067 => x"38b5a408",
  1068 => x"fe06b5a4",
  1069 => x"0c800bb5",
  1070 => x"ac0cba88",
  1071 => x"519cf72d",
  1072 => x"b3fc0855",
  1073 => x"b3fc08ff",
  1074 => x"24fdea38",
  1075 => x"76802e94",
  1076 => x"3881ed52",
  1077 => x"ba88519e",
  1078 => x"d62db5a8",
  1079 => x"0852ba88",
  1080 => x"519ed62d",
  1081 => x"805372b3",
  1082 => x"fc0c029c",
  1083 => x"050d0402",
  1084 => x"fc050d80",
  1085 => x"51800ba9",
  1086 => x"fc1281b7",
  1087 => x"2d811151",
  1088 => x"81ff7125",
  1089 => x"f0380284",
  1090 => x"050d0402",
  1091 => x"f4050d74",
  1092 => x"51a2c82d",
  1093 => x"a9fc1180",
  1094 => x"f52d7081",
  1095 => x"ff0671fd",
  1096 => x"06525452",
  1097 => x"71a9fc12",
  1098 => x"81b72da2",
  1099 => x"c22d72b3",
  1100 => x"fc0c028c",
  1101 => x"050d0471",
  1102 => x"980c04ff",
  1103 => x"b008b3fc",
  1104 => x"0c04810b",
  1105 => x"ffb00c04",
  1106 => x"800bffb0",
  1107 => x"0c0402e8",
  1108 => x"050d7878",
  1109 => x"71545753",
  1110 => x"72802584",
  1111 => x"38831352",
  1112 => x"71822cff",
  1113 => x"055372ff",
  1114 => x"2e80c038",
  1115 => x"75708405",
  1116 => x"57085487",
  1117 => x"55739c2a",
  1118 => x"b00552b9",
  1119 => x"72278438",
  1120 => x"87125271",
  1121 => x"5195c92d",
  1122 => x"73842bff",
  1123 => x"16565474",
  1124 => x"8025e238",
  1125 => x"a05195c9",
  1126 => x"2d728706",
  1127 => x"52718638",
  1128 => x"8a5195c9",
  1129 => x"2dff1353",
  1130 => x"a2e6048a",
  1131 => x"5195c92d",
  1132 => x"0298050d",
  1133 => x"04b48808",
  1134 => x"02b4880c",
  1135 => x"ff3d0d80",
  1136 => x"0bb48808",
  1137 => x"fc050cb4",
  1138 => x"88088805",
  1139 => x"088106ff",
  1140 => x"11700970",
  1141 => x"b488088c",
  1142 => x"050806b4",
  1143 => x"8808fc05",
  1144 => x"0811b488",
  1145 => x"08fc050c",
  1146 => x"b4880888",
  1147 => x"0508812a",
  1148 => x"b4880888",
  1149 => x"050cb488",
  1150 => x"088c0508",
  1151 => x"10b48808",
  1152 => x"8c050c51",
  1153 => x"515151b4",
  1154 => x"88088805",
  1155 => x"08802e84",
  1156 => x"38ffb439",
  1157 => x"b48808fc",
  1158 => x"050870b3",
  1159 => x"fc0c5183",
  1160 => x"3d0db488",
  1161 => x"0c040000",
  1162 => x"00ffffff",
  1163 => x"ff00ffff",
  1164 => x"ffff00ff",
  1165 => x"ffffff00",
  1166 => x"496e6974",
  1167 => x"69616c69",
  1168 => x"73696e67",
  1169 => x"2050532f",
  1170 => x"3220696e",
  1171 => x"74657266",
  1172 => x"6163652e",
  1173 => x"2e2e0a00",
  1174 => x"496e6974",
  1175 => x"69616c69",
  1176 => x"7a696e67",
  1177 => x"20534420",
  1178 => x"63617264",
  1179 => x"0a000000",
  1180 => x"48756e74",
  1181 => x"696e6720",
  1182 => x"666f7220",
  1183 => x"70617274",
  1184 => x"6974696f",
  1185 => x"6e0a0000",
  1186 => x"42494f53",
  1187 => x"5041434b",
  1188 => x"524f4d00",
  1189 => x"4f70656e",
  1190 => x"65642066",
  1191 => x"696c652c",
  1192 => x"206c6f61",
  1193 => x"64696e67",
  1194 => x"2e2e2e0a",
  1195 => x"00000000",
  1196 => x"52656164",
  1197 => x"20626c6f",
  1198 => x"636b2066",
  1199 => x"61696c65",
  1200 => x"640a0000",
  1201 => x"4c6f6164",
  1202 => x"696e6720",
  1203 => x"42494f53",
  1204 => x"20666169",
  1205 => x"6c65640a",
  1206 => x"00000000",
  1207 => x"52656164",
  1208 => x"696e6720",
  1209 => x"4d42520a",
  1210 => x"00000000",
  1211 => x"52656164",
  1212 => x"206f6620",
  1213 => x"4d425220",
  1214 => x"6661696c",
  1215 => x"65640a00",
  1216 => x"4d425220",
  1217 => x"73756363",
  1218 => x"65737366",
  1219 => x"756c6c79",
  1220 => x"20726561",
  1221 => x"640a0000",
  1222 => x"46415431",
  1223 => x"36202020",
  1224 => x"00000000",
  1225 => x"46415433",
  1226 => x"32202020",
  1227 => x"00000000",
  1228 => x"50617274",
  1229 => x"6974696f",
  1230 => x"6e636f75",
  1231 => x"6e742025",
  1232 => x"640a0000",
  1233 => x"4e6f2070",
  1234 => x"61727469",
  1235 => x"74696f6e",
  1236 => x"20736967",
  1237 => x"6e617475",
  1238 => x"72652066",
  1239 => x"6f756e64",
  1240 => x"0a000000",
  1241 => x"52656164",
  1242 => x"696e6720",
  1243 => x"626f6f74",
  1244 => x"20736563",
  1245 => x"746f7220",
  1246 => x"25640a00",
  1247 => x"52656164",
  1248 => x"20626f6f",
  1249 => x"74207365",
  1250 => x"63746f72",
  1251 => x"2066726f",
  1252 => x"6d206669",
  1253 => x"72737420",
  1254 => x"70617274",
  1255 => x"6974696f",
  1256 => x"6e0a0000",
  1257 => x"48756e74",
  1258 => x"696e6720",
  1259 => x"666f7220",
  1260 => x"66696c65",
  1261 => x"73797374",
  1262 => x"656d0a00",
  1263 => x"556e7375",
  1264 => x"70706f72",
  1265 => x"74656420",
  1266 => x"70617274",
  1267 => x"6974696f",
  1268 => x"6e207479",
  1269 => x"7065210d",
  1270 => x"00000000",
  1271 => x"436c7573",
  1272 => x"74657220",
  1273 => x"73697a65",
  1274 => x"3a202564",
  1275 => x"2c20436c",
  1276 => x"75737465",
  1277 => x"72206d61",
  1278 => x"736b2c20",
  1279 => x"25640a00",
  1280 => x"47657443",
  1281 => x"6c757374",
  1282 => x"65722072",
  1283 => x"65616469",
  1284 => x"6e672073",
  1285 => x"6563746f",
  1286 => x"72202564",
  1287 => x"0a000000",
  1288 => x"52656164",
  1289 => x"696e6720",
  1290 => x"64697265",
  1291 => x"63746f72",
  1292 => x"79207365",
  1293 => x"63746f72",
  1294 => x"2025640a",
  1295 => x"00000000",
  1296 => x"47657446",
  1297 => x"41544c69",
  1298 => x"6e6b2072",
  1299 => x"65747572",
  1300 => x"6e656420",
  1301 => x"25640a00",
  1302 => x"436d645f",
  1303 => x"696e6974",
  1304 => x"0a000000",
  1305 => x"636d645f",
  1306 => x"434d4438",
  1307 => x"20726573",
  1308 => x"706f6e73",
  1309 => x"653a2025",
  1310 => x"640a0000",
  1311 => x"434d4438",
  1312 => x"5f342072",
  1313 => x"6573706f",
  1314 => x"6e73653a",
  1315 => x"2025640a",
  1316 => x"00000000",
  1317 => x"53444843",
  1318 => x"20496e69",
  1319 => x"7469616c",
  1320 => x"697a6174",
  1321 => x"696f6e20",
  1322 => x"6572726f",
  1323 => x"72210a00",
  1324 => x"434d4435",
  1325 => x"38202564",
  1326 => x"0a202000",
  1327 => x"434d4435",
  1328 => x"385f3220",
  1329 => x"25640a20",
  1330 => x"20000000",
  1331 => x"53504920",
  1332 => x"496e6974",
  1333 => x"28290a00",
  1334 => x"52656164",
  1335 => x"20636f6d",
  1336 => x"6d616e64",
  1337 => x"20666169",
  1338 => x"6c656420",
  1339 => x"61742025",
  1340 => x"64202825",
  1341 => x"64290a00",
  1342 => x"ffffe000",
  1343 => x"00000000",
  1344 => x"00000000",
  1345 => x"00000000",
  1346 => x"00000000",
  1347 => x"00000000",
  1348 => x"00000000",
  1349 => x"00000000",
  1350 => x"00000000",
  1351 => x"00000000",
  1352 => x"00000000",
  1353 => x"00000000",
  1354 => x"00000000",
  1355 => x"00000000",
  1356 => x"00000000",
  1357 => x"00000000",
  1358 => x"00000000",
  1359 => x"00000000",
  1360 => x"00000000",
  1361 => x"00000000",
  1362 => x"00000000",
  1363 => x"00000000",
  1364 => x"00000000",
  1365 => x"00000000",
  1366 => x"00000000",
  1367 => x"00000000",
  1368 => x"00000000",
  1369 => x"00000000",
  1370 => x"00000000",
  1371 => x"00000000",
  1372 => x"00000000",
  1373 => x"00000000",
  1374 => x"00000000",
  1375 => x"00000000",
  1376 => x"00000000",
  1377 => x"00000000",
  1378 => x"00000000",
  1379 => x"00000000",
  1380 => x"00000000",
  1381 => x"00000000",
  1382 => x"00000000",
  1383 => x"00000000",
  1384 => x"00000000",
  1385 => x"00000000",
  1386 => x"00000000",
  1387 => x"00000000",
  1388 => x"00000000",
  1389 => x"00000000",
  1390 => x"00000000",
  1391 => x"00000000",
  1392 => x"00000000",
  1393 => x"00000000",
  1394 => x"00000000",
  1395 => x"00000000",
  1396 => x"00000000",
  1397 => x"00000000",
  1398 => x"00000000",
  1399 => x"00000000",
  1400 => x"00000000",
  1401 => x"00000000",
  1402 => x"00000000",
  1403 => x"00000000",
  1404 => x"00000000",
  1405 => x"00000000",
  1406 => x"00000000",
  1407 => x"00000000",
  1408 => x"00000000",
  1409 => x"00000000",
  1410 => x"00000000",
  1411 => x"00000000",
  1412 => x"00000000",
  1413 => x"00000000",
  1414 => x"00000000",
  1415 => x"00000000",
  1416 => x"00000000",
  1417 => x"00000000",
  1418 => x"00000000",
  1419 => x"00000000",
  1420 => x"00000009",
  1421 => x"00000000",
  1422 => x"00000000",
  1423 => x"00000000",
  1424 => x"00000000",
  1425 => x"00000000",
  1426 => x"00000000",
  1427 => x"00000000",
  1428 => x"00000071",
  1429 => x"00000031",
  1430 => x"00000000",
  1431 => x"00000000",
  1432 => x"00000000",
  1433 => x"0000007a",
  1434 => x"00000073",
  1435 => x"00000061",
  1436 => x"00000077",
  1437 => x"00000032",
  1438 => x"00000000",
  1439 => x"00000000",
  1440 => x"00000063",
  1441 => x"00000078",
  1442 => x"00000064",
  1443 => x"00000065",
  1444 => x"00000034",
  1445 => x"00000033",
  1446 => x"00000000",
  1447 => x"00000000",
  1448 => x"00000020",
  1449 => x"00000076",
  1450 => x"00000066",
  1451 => x"00000074",
  1452 => x"00000072",
  1453 => x"00000035",
  1454 => x"00000000",
  1455 => x"00000000",
  1456 => x"0000006e",
  1457 => x"00000062",
  1458 => x"00000068",
  1459 => x"00000067",
  1460 => x"00000079",
  1461 => x"00000036",
  1462 => x"00000000",
  1463 => x"00000000",
  1464 => x"00000000",
  1465 => x"0000006d",
  1466 => x"0000006a",
  1467 => x"00000075",
  1468 => x"00000037",
  1469 => x"00000038",
  1470 => x"00000000",
  1471 => x"00000000",
  1472 => x"0000002c",
  1473 => x"0000006b",
  1474 => x"00000069",
  1475 => x"0000006f",
  1476 => x"00000030",
  1477 => x"00000039",
  1478 => x"00000000",
  1479 => x"00000000",
  1480 => x"0000002e",
  1481 => x"0000002f",
  1482 => x"0000006c",
  1483 => x"0000003b",
  1484 => x"00000070",
  1485 => x"0000002d",
  1486 => x"00000000",
  1487 => x"00000000",
  1488 => x"00000000",
  1489 => x"00000027",
  1490 => x"00000000",
  1491 => x"0000005b",
  1492 => x"0000003d",
  1493 => x"00000000",
  1494 => x"00000000",
  1495 => x"00000000",
  1496 => x"00000000",
  1497 => x"0000000a",
  1498 => x"0000005d",
  1499 => x"00000000",
  1500 => x"00000023",
  1501 => x"00000000",
  1502 => x"00000000",
  1503 => x"00000000",
  1504 => x"00000000",
  1505 => x"00000000",
  1506 => x"00000000",
  1507 => x"00000000",
  1508 => x"00000000",
  1509 => x"00000008",
  1510 => x"00000000",
  1511 => x"00000000",
  1512 => x"00000031",
  1513 => x"00000000",
  1514 => x"00000034",
  1515 => x"00000037",
  1516 => x"00000000",
  1517 => x"00000000",
  1518 => x"00000000",
  1519 => x"00000030",
  1520 => x"0000002e",
  1521 => x"00000032",
  1522 => x"00000035",
  1523 => x"00000036",
  1524 => x"00000038",
  1525 => x"0000001b",
  1526 => x"00000000",
  1527 => x"00000000",
  1528 => x"0000002b",
  1529 => x"00000033",
  1530 => x"00000000",
  1531 => x"0000002a",
  1532 => x"00000039",
  1533 => x"00000000",
  1534 => x"00000000",
  1535 => x"00000000",
  1536 => x"00000000",
  1537 => x"00000000",
  1538 => x"00000000",
  1539 => x"00000000",
  1540 => x"00000000",
  1541 => x"00000000",
  1542 => x"00000000",
  1543 => x"00000000",
  1544 => x"00000000",
  1545 => x"00000000",
  1546 => x"00000000",
  1547 => x"00000000",
  1548 => x"00000008",
  1549 => x"00000000",
  1550 => x"00000000",
  1551 => x"00000000",
  1552 => x"00000000",
  1553 => x"00000000",
  1554 => x"00000000",
  1555 => x"00000000",
  1556 => x"00000051",
  1557 => x"00000021",
  1558 => x"00000000",
  1559 => x"00000000",
  1560 => x"00000000",
  1561 => x"0000005a",
  1562 => x"00000053",
  1563 => x"00000041",
  1564 => x"00000057",
  1565 => x"00000022",
  1566 => x"00000000",
  1567 => x"00000000",
  1568 => x"00000043",
  1569 => x"00000058",
  1570 => x"00000044",
  1571 => x"00000045",
  1572 => x"00000024",
  1573 => x"000000a3",
  1574 => x"00000000",
  1575 => x"00000000",
  1576 => x"00000020",
  1577 => x"00000056",
  1578 => x"00000046",
  1579 => x"00000054",
  1580 => x"00000052",
  1581 => x"00000025",
  1582 => x"00000000",
  1583 => x"00000000",
  1584 => x"0000004e",
  1585 => x"00000042",
  1586 => x"00000048",
  1587 => x"00000047",
  1588 => x"00000059",
  1589 => x"0000005e",
  1590 => x"00000000",
  1591 => x"00000000",
  1592 => x"00000000",
  1593 => x"0000004d",
  1594 => x"0000004a",
  1595 => x"00000055",
  1596 => x"00000026",
  1597 => x"0000002a",
  1598 => x"00000000",
  1599 => x"00000000",
  1600 => x"0000003c",
  1601 => x"0000004b",
  1602 => x"00000049",
  1603 => x"0000004f",
  1604 => x"00000029",
  1605 => x"00000028",
  1606 => x"00000000",
  1607 => x"00000000",
  1608 => x"0000003e",
  1609 => x"0000003f",
  1610 => x"0000004c",
  1611 => x"0000003a",
  1612 => x"00000050",
  1613 => x"0000005f",
  1614 => x"00000000",
  1615 => x"00000000",
  1616 => x"00000000",
  1617 => x"0000003f",
  1618 => x"00000000",
  1619 => x"0000007b",
  1620 => x"0000002b",
  1621 => x"00000000",
  1622 => x"00000000",
  1623 => x"00000000",
  1624 => x"00000000",
  1625 => x"0000000a",
  1626 => x"0000007d",
  1627 => x"00000000",
  1628 => x"0000007e",
  1629 => x"00000000",
  1630 => x"00000000",
  1631 => x"00000000",
  1632 => x"00000000",
  1633 => x"00000000",
  1634 => x"00000000",
  1635 => x"00000000",
  1636 => x"00000000",
  1637 => x"00000009",
  1638 => x"00000000",
  1639 => x"00000000",
  1640 => x"00000031",
  1641 => x"00000000",
  1642 => x"00000034",
  1643 => x"00000037",
  1644 => x"00000000",
  1645 => x"00000000",
  1646 => x"00000000",
  1647 => x"00000030",
  1648 => x"0000002e",
  1649 => x"00000032",
  1650 => x"00000035",
  1651 => x"00000036",
  1652 => x"00000038",
  1653 => x"0000001b",
  1654 => x"00000000",
  1655 => x"00000000",
  1656 => x"0000002b",
  1657 => x"00000033",
  1658 => x"00000000",
  1659 => x"0000002a",
  1660 => x"00000039",
  1661 => x"00000000",
  1662 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

