-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b0bb1",
     9 => x"d8080b0b",
    10 => x"0bb1dc08",
    11 => x"0b0b0bb1",
    12 => x"e0080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"b1e00c0b",
    16 => x"0b0bb1dc",
    17 => x"0c0b0b0b",
    18 => x"b1d80c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0ba8b4",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"b1d870b7",
    57 => x"b4278b38",
    58 => x"80717084",
    59 => x"05530c81",
    60 => x"e2048c51",
    61 => x"8af80402",
    62 => x"fc050df8",
    63 => x"80518f0b",
    64 => x"b1e80c9f",
    65 => x"0bb1ec0c",
    66 => x"a0717081",
    67 => x"055334b1",
    68 => x"ec08ff05",
    69 => x"b1ec0cb1",
    70 => x"ec088025",
    71 => x"eb38b1e8",
    72 => x"08ff05b1",
    73 => x"e80cb1e8",
    74 => x"088025d7",
    75 => x"38028405",
    76 => x"0d0402f0",
    77 => x"050df880",
    78 => x"53f8a054",
    79 => x"83bf5273",
    80 => x"70810555",
    81 => x"33517073",
    82 => x"70810555",
    83 => x"34ff1252",
    84 => x"718025eb",
    85 => x"38fbc053",
    86 => x"9f52a073",
    87 => x"70810555",
    88 => x"34ff1252",
    89 => x"718025f2",
    90 => x"38029005",
    91 => x"0d0402f4",
    92 => x"050d7453",
    93 => x"8e0bb1e8",
    94 => x"08258f38",
    95 => x"82b22db1",
    96 => x"e808ff05",
    97 => x"b1e80c82",
    98 => x"f404b1e8",
    99 => x"08b1ec08",
   100 => x"5351728a",
   101 => x"2e098106",
   102 => x"b7387151",
   103 => x"719f24a0",
   104 => x"38b1e808",
   105 => x"a02911f8",
   106 => x"80115151",
   107 => x"a07134b1",
   108 => x"ec088105",
   109 => x"b1ec0cb1",
   110 => x"ec08519f",
   111 => x"7125e238",
   112 => x"800bb1ec",
   113 => x"0cb1e808",
   114 => x"8105b1e8",
   115 => x"0c83e404",
   116 => x"70a02912",
   117 => x"f8801151",
   118 => x"51727134",
   119 => x"b1ec0881",
   120 => x"05b1ec0c",
   121 => x"b1ec08a0",
   122 => x"2e098106",
   123 => x"8e38800b",
   124 => x"b1ec0cb1",
   125 => x"e8088105",
   126 => x"b1e80c02",
   127 => x"8c050d04",
   128 => x"02e8050d",
   129 => x"77795656",
   130 => x"880bfc16",
   131 => x"77712c8f",
   132 => x"06545254",
   133 => x"80537272",
   134 => x"25953871",
   135 => x"53fbe014",
   136 => x"51877134",
   137 => x"8114ff14",
   138 => x"545472f1",
   139 => x"387153f9",
   140 => x"1576712c",
   141 => x"87065351",
   142 => x"71802e8b",
   143 => x"38fbe014",
   144 => x"51717134",
   145 => x"81145472",
   146 => x"8e249538",
   147 => x"8f733153",
   148 => x"fbe01451",
   149 => x"a0713481",
   150 => x"14ff1454",
   151 => x"5472f138",
   152 => x"0298050d",
   153 => x"0402ec05",
   154 => x"0d800bb1",
   155 => x"f00cf68c",
   156 => x"08f69008",
   157 => x"71882c56",
   158 => x"5481ff06",
   159 => x"52737225",
   160 => x"88387154",
   161 => x"820bb1f0",
   162 => x"0c72882c",
   163 => x"7381ff06",
   164 => x"54557473",
   165 => x"258b3872",
   166 => x"b1f00884",
   167 => x"07b1f00c",
   168 => x"550b0b0b",
   169 => x"afbc0882",
   170 => x"0574712b",
   171 => x"86a07125",
   172 => x"83713170",
   173 => x"0b0b0baf",
   174 => x"bc0c8171",
   175 => x"2bff05f6",
   176 => x"880cfecc",
   177 => x"13ff122c",
   178 => x"798829ff",
   179 => x"94057081",
   180 => x"2cb1f008",
   181 => x"52595256",
   182 => x"51525551",
   183 => x"76802e85",
   184 => x"38708107",
   185 => x"5170f694",
   186 => x"0c710981",
   187 => x"05f6800c",
   188 => x"72098105",
   189 => x"f6840c02",
   190 => x"94050d04",
   191 => x"02f4050d",
   192 => x"74537270",
   193 => x"81055480",
   194 => x"f52d5271",
   195 => x"802e8938",
   196 => x"715182ee",
   197 => x"2d868204",
   198 => x"028c050d",
   199 => x"0402f805",
   200 => x"0da28d2d",
   201 => x"80da51a3",
   202 => x"c42db1d8",
   203 => x"08812a70",
   204 => x"81065152",
   205 => x"71802ee9",
   206 => x"38028805",
   207 => x"0d0402f4",
   208 => x"050db7a4",
   209 => x"0881c406",
   210 => x"b0c00b80",
   211 => x"f52d5252",
   212 => x"70802e86",
   213 => x"38718480",
   214 => x"0752aff8",
   215 => x"0b80f52d",
   216 => x"7207b090",
   217 => x"0b80f52d",
   218 => x"70812a70",
   219 => x"81065153",
   220 => x"54527080",
   221 => x"2e863871",
   222 => x"82800752",
   223 => x"72810651",
   224 => x"70802e85",
   225 => x"38718807",
   226 => x"52b09c0b",
   227 => x"80f52d70",
   228 => x"842b7307",
   229 => x"8432b1d8",
   230 => x"0c51028c",
   231 => x"050d0402",
   232 => x"f4050d74",
   233 => x"708432b7",
   234 => x"a40c7083",
   235 => x"06525370",
   236 => x"aff00b88",
   237 => x"0581b72d",
   238 => x"72892a70",
   239 => x"81065151",
   240 => x"70b0c00b",
   241 => x"81b72d72",
   242 => x"832a8106",
   243 => x"73882a70",
   244 => x"81065152",
   245 => x"5270802e",
   246 => x"85387182",
   247 => x"075271b0",
   248 => x"900b81b7",
   249 => x"2d72842c",
   250 => x"70830651",
   251 => x"5170b09c",
   252 => x"0b81b72d",
   253 => x"70b1d80c",
   254 => x"028c050d",
   255 => x"0402d405",
   256 => x"0dab8051",
   257 => x"85fc2d9a",
   258 => x"8e2db1d8",
   259 => x"08802e82",
   260 => x"ab3886be",
   261 => x"2db1d808",
   262 => x"538ce92d",
   263 => x"b1d80854",
   264 => x"b1d80880",
   265 => x"2e829738",
   266 => x"9cd12db1",
   267 => x"d808802e",
   268 => x"8738ab98",
   269 => x"5188c504",
   270 => x"95f02db1",
   271 => x"d808802e",
   272 => x"9c38abd8",
   273 => x"5185fc2d",
   274 => x"869d2d72",
   275 => x"84075381",
   276 => x"0bfec40c",
   277 => x"72fec00c",
   278 => x"7251879f",
   279 => x"2d840bfe",
   280 => x"c40caca0",
   281 => x"5185fc2d",
   282 => x"acb852b1",
   283 => x"f8519385",
   284 => x"2db1d808",
   285 => x"9838acc4",
   286 => x"5185fc2d",
   287 => x"acdc52b1",
   288 => x"f8519385",
   289 => x"2db1d808",
   290 => x"802e81b0",
   291 => x"38ace851",
   292 => x"85fc2db1",
   293 => x"fc085780",
   294 => x"77595a76",
   295 => x"7a2e8b38",
   296 => x"811a7881",
   297 => x"2a595a77",
   298 => x"f738f71a",
   299 => x"5a807725",
   300 => x"81803879",
   301 => x"52775184",
   302 => x"802db284",
   303 => x"52b1f851",
   304 => x"95ca2db1",
   305 => x"d80853b1",
   306 => x"d808802e",
   307 => x"80c938b2",
   308 => x"845b8059",
   309 => x"8a84047a",
   310 => x"7084055c",
   311 => x"087081ff",
   312 => x"0671882c",
   313 => x"7081ff06",
   314 => x"73902c70",
   315 => x"81ff0675",
   316 => x"982afec8",
   317 => x"0cfec80c",
   318 => x"58fec80c",
   319 => x"57fec80c",
   320 => x"841a5a53",
   321 => x"76538480",
   322 => x"77258438",
   323 => x"84805372",
   324 => x"7924c438",
   325 => x"8aa204ad",
   326 => x"845185fc",
   327 => x"2d72548a",
   328 => x"be04b1f8",
   329 => x"51959d2d",
   330 => x"fc801781",
   331 => x"19595789",
   332 => x"ad04820b",
   333 => x"fec40c81",
   334 => x"548abe04",
   335 => x"805473b1",
   336 => x"d80c02ac",
   337 => x"050d0402",
   338 => x"f8050da4",
   339 => x"942d81f7",
   340 => x"2d815184",
   341 => x"e52dfec4",
   342 => x"5281720c",
   343 => x"a1da2da1",
   344 => x"da2d8472",
   345 => x"0c87fd2d",
   346 => x"afc051a5",
   347 => x"ad2d8051",
   348 => x"84e52d02",
   349 => x"88050d04",
   350 => x"02f4050d",
   351 => x"84b95187",
   352 => x"9f2d810b",
   353 => x"fec40c84",
   354 => x"b90bfec0",
   355 => x"0c840bfe",
   356 => x"c40ca1f5",
   357 => x"2da4882d",
   358 => x"a1da2da1",
   359 => x"da2d81f7",
   360 => x"2d815184",
   361 => x"e52da1da",
   362 => x"2da1da2d",
   363 => x"815184e5",
   364 => x"2d87fd2d",
   365 => x"b1d80880",
   366 => x"2e80db38",
   367 => x"805184e5",
   368 => x"2dafc051",
   369 => x"a5ad2da2",
   370 => x"8d2da5bd",
   371 => x"2db1d808",
   372 => x"5386be2d",
   373 => x"b1d808fe",
   374 => x"c00c86be",
   375 => x"2db1d808",
   376 => x"b1f4082e",
   377 => x"9c38b1d8",
   378 => x"08b1f40c",
   379 => x"85527251",
   380 => x"84e52da1",
   381 => x"da2da1da",
   382 => x"2dff1252",
   383 => x"718025ee",
   384 => x"3872802e",
   385 => x"89388a0b",
   386 => x"fec40c8b",
   387 => x"c704820b",
   388 => x"fec40c8b",
   389 => x"c704ad98",
   390 => x"5185fc2d",
   391 => x"820bfec4",
   392 => x"0c800bb1",
   393 => x"d80c028c",
   394 => x"050d0402",
   395 => x"e8050d77",
   396 => x"797b5855",
   397 => x"55805372",
   398 => x"7625a338",
   399 => x"74708105",
   400 => x"5680f52d",
   401 => x"74708105",
   402 => x"5680f52d",
   403 => x"52527171",
   404 => x"2e863881",
   405 => x"518ce004",
   406 => x"8113538c",
   407 => x"b7048051",
   408 => x"70b1d80c",
   409 => x"0298050d",
   410 => x"0402d805",
   411 => x"0d800bb6",
   412 => x"8c0cb284",
   413 => x"5280519b",
   414 => x"ae2db1d8",
   415 => x"0854b1d8",
   416 => x"088c38ad",
   417 => x"b05185fc",
   418 => x"2d735592",
   419 => x"8e048056",
   420 => x"810bb6b0",
   421 => x"0c8853ad",
   422 => x"c452b2ba",
   423 => x"518cab2d",
   424 => x"b1d80876",
   425 => x"2e098106",
   426 => x"8738b1d8",
   427 => x"08b6b00c",
   428 => x"8853add0",
   429 => x"52b2d651",
   430 => x"8cab2db1",
   431 => x"d8088738",
   432 => x"b1d808b6",
   433 => x"b00cb6b0",
   434 => x"0852addc",
   435 => x"519ecb2d",
   436 => x"b6b00880",
   437 => x"2e80f638",
   438 => x"b5ca0b80",
   439 => x"f52db5cb",
   440 => x"0b80f52d",
   441 => x"71982b71",
   442 => x"902b07b5",
   443 => x"cc0b80f5",
   444 => x"2d70882b",
   445 => x"7207b5cd",
   446 => x"0b80f52d",
   447 => x"7107b682",
   448 => x"0b80f52d",
   449 => x"b6830b80",
   450 => x"f52d7188",
   451 => x"2b07535f",
   452 => x"54525a56",
   453 => x"57557381",
   454 => x"abaa2e09",
   455 => x"81068d38",
   456 => x"75519da0",
   457 => x"2db1d808",
   458 => x"568eb904",
   459 => x"7382d4d5",
   460 => x"2e8738ad",
   461 => x"f4518efa",
   462 => x"04b28452",
   463 => x"75519bae",
   464 => x"2db1d808",
   465 => x"55b1d808",
   466 => x"802e83c2",
   467 => x"388853ad",
   468 => x"d052b2d6",
   469 => x"518cab2d",
   470 => x"b1d80889",
   471 => x"38810bb6",
   472 => x"8c0c8f80",
   473 => x"048853ad",
   474 => x"c452b2ba",
   475 => x"518cab2d",
   476 => x"b1d80880",
   477 => x"2e8a38ae",
   478 => x"945185fc",
   479 => x"2d8fda04",
   480 => x"b6820b80",
   481 => x"f52d5473",
   482 => x"80d52e09",
   483 => x"810680ca",
   484 => x"38b6830b",
   485 => x"80f52d54",
   486 => x"7381aa2e",
   487 => x"098106ba",
   488 => x"38800bb2",
   489 => x"840b80f5",
   490 => x"2d565474",
   491 => x"81e92e83",
   492 => x"38815474",
   493 => x"81eb2e8c",
   494 => x"38805573",
   495 => x"752e0981",
   496 => x"0682cb38",
   497 => x"b28f0b80",
   498 => x"f52d5574",
   499 => x"8d38b290",
   500 => x"0b80f52d",
   501 => x"5473822e",
   502 => x"86388055",
   503 => x"928e04b2",
   504 => x"910b80f5",
   505 => x"2d70b684",
   506 => x"0cff05b6",
   507 => x"880cb292",
   508 => x"0b80f52d",
   509 => x"b2930b80",
   510 => x"f52d5876",
   511 => x"05778280",
   512 => x"290570b6",
   513 => x"900cb294",
   514 => x"0b80f52d",
   515 => x"70b6a40c",
   516 => x"b68c0859",
   517 => x"57587680",
   518 => x"2e81a338",
   519 => x"8853add0",
   520 => x"52b2d651",
   521 => x"8cab2db1",
   522 => x"d80881e2",
   523 => x"38b68408",
   524 => x"70842bb6",
   525 => x"a80c70b6",
   526 => x"a00cb2a9",
   527 => x"0b80f52d",
   528 => x"b2a80b80",
   529 => x"f52d7182",
   530 => x"802905b2",
   531 => x"aa0b80f5",
   532 => x"2d708480",
   533 => x"802912b2",
   534 => x"ab0b80f5",
   535 => x"2d708180",
   536 => x"0a291270",
   537 => x"b6ac0cb6",
   538 => x"a4087129",
   539 => x"b6900805",
   540 => x"70b6940c",
   541 => x"b2b10b80",
   542 => x"f52db2b0",
   543 => x"0b80f52d",
   544 => x"71828029",
   545 => x"05b2b20b",
   546 => x"80f52d70",
   547 => x"84808029",
   548 => x"12b2b30b",
   549 => x"80f52d70",
   550 => x"982b81f0",
   551 => x"0a067205",
   552 => x"70b6980c",
   553 => x"fe117e29",
   554 => x"7705b69c",
   555 => x"0c525952",
   556 => x"43545e51",
   557 => x"5259525d",
   558 => x"57595792",
   559 => x"8c04b296",
   560 => x"0b80f52d",
   561 => x"b2950b80",
   562 => x"f52d7182",
   563 => x"80290570",
   564 => x"b6a80c70",
   565 => x"a02983ff",
   566 => x"0570892a",
   567 => x"70b6a00c",
   568 => x"b29b0b80",
   569 => x"f52db29a",
   570 => x"0b80f52d",
   571 => x"71828029",
   572 => x"0570b6ac",
   573 => x"0c7b7129",
   574 => x"1e70b69c",
   575 => x"0c7db698",
   576 => x"0c7305b6",
   577 => x"940c555e",
   578 => x"51515555",
   579 => x"815574b1",
   580 => x"d80c02a8",
   581 => x"050d0402",
   582 => x"ec050d76",
   583 => x"70872c71",
   584 => x"80ff0655",
   585 => x"5654b68c",
   586 => x"088a3873",
   587 => x"882c7481",
   588 => x"ff065455",
   589 => x"b28452b6",
   590 => x"90081551",
   591 => x"9bae2db1",
   592 => x"d80854b1",
   593 => x"d808802e",
   594 => x"b338b68c",
   595 => x"08802e98",
   596 => x"38728429",
   597 => x"b2840570",
   598 => x"0852539d",
   599 => x"a02db1d8",
   600 => x"08f00a06",
   601 => x"5392fa04",
   602 => x"7210b284",
   603 => x"057080e0",
   604 => x"2d52539d",
   605 => x"d02db1d8",
   606 => x"08537254",
   607 => x"73b1d80c",
   608 => x"0294050d",
   609 => x"0402c805",
   610 => x"0d7f615f",
   611 => x"5b800bb6",
   612 => x"9808b69c",
   613 => x"08595d56",
   614 => x"b68c0876",
   615 => x"2e8a38b6",
   616 => x"8408842b",
   617 => x"5893ae04",
   618 => x"b6a00884",
   619 => x"2b588059",
   620 => x"78782781",
   621 => x"a938788f",
   622 => x"06a01757",
   623 => x"54738f38",
   624 => x"b2845276",
   625 => x"51811757",
   626 => x"9bae2db2",
   627 => x"84568076",
   628 => x"80f52d56",
   629 => x"5474742e",
   630 => x"83388154",
   631 => x"7481e52e",
   632 => x"80f63881",
   633 => x"70750655",
   634 => x"5d73802e",
   635 => x"80ea388b",
   636 => x"1680f52d",
   637 => x"98065a79",
   638 => x"80de388b",
   639 => x"537d5275",
   640 => x"518cab2d",
   641 => x"b1d80880",
   642 => x"cf389c16",
   643 => x"08519da0",
   644 => x"2db1d808",
   645 => x"841c0c9a",
   646 => x"1680e02d",
   647 => x"519dd02d",
   648 => x"b1d808b1",
   649 => x"d808881d",
   650 => x"0cb1d808",
   651 => x"5555b68c",
   652 => x"08802e98",
   653 => x"38941680",
   654 => x"e02d519d",
   655 => x"d02db1d8",
   656 => x"08902b83",
   657 => x"fff00a06",
   658 => x"70165154",
   659 => x"73881c0c",
   660 => x"797b0c7c",
   661 => x"54959404",
   662 => x"81195993",
   663 => x"b004b68c",
   664 => x"08802eae",
   665 => x"387b5192",
   666 => x"972db1d8",
   667 => x"08b1d808",
   668 => x"80ffffff",
   669 => x"f806555c",
   670 => x"7380ffff",
   671 => x"fff82e92",
   672 => x"38b1d808",
   673 => x"fe05b684",
   674 => x"0829b694",
   675 => x"08055793",
   676 => x"ae048054",
   677 => x"73b1d80c",
   678 => x"02b8050d",
   679 => x"0402f405",
   680 => x"0d747008",
   681 => x"8105710c",
   682 => x"7008b688",
   683 => x"08065353",
   684 => x"718e3888",
   685 => x"13085192",
   686 => x"972db1d8",
   687 => x"0888140c",
   688 => x"810bb1d8",
   689 => x"0c028c05",
   690 => x"0d0402f0",
   691 => x"050d7588",
   692 => x"1108fe05",
   693 => x"b6840829",
   694 => x"b6940811",
   695 => x"7208b688",
   696 => x"08060579",
   697 => x"55535454",
   698 => x"9bae2d02",
   699 => x"90050d04",
   700 => x"b68c08b1",
   701 => x"d80c0402",
   702 => x"f4050dd4",
   703 => x"5281ff72",
   704 => x"0c710853",
   705 => x"81ff720c",
   706 => x"72882b83",
   707 => x"fe800672",
   708 => x"087081ff",
   709 => x"06515253",
   710 => x"81ff720c",
   711 => x"72710788",
   712 => x"2b720870",
   713 => x"81ff0651",
   714 => x"525381ff",
   715 => x"720c7271",
   716 => x"07882b72",
   717 => x"087081ff",
   718 => x"067207b1",
   719 => x"d80c5253",
   720 => x"028c050d",
   721 => x"0402f405",
   722 => x"0d747671",
   723 => x"81ff06d4",
   724 => x"0c5353b6",
   725 => x"b4088538",
   726 => x"71892b52",
   727 => x"71982ad4",
   728 => x"0c71902a",
   729 => x"7081ff06",
   730 => x"d40c5171",
   731 => x"882a7081",
   732 => x"ff06d40c",
   733 => x"517181ff",
   734 => x"06d40c72",
   735 => x"902a7081",
   736 => x"ff06d40c",
   737 => x"51d40870",
   738 => x"81ff0651",
   739 => x"5182b8bf",
   740 => x"527081ff",
   741 => x"2e098106",
   742 => x"943881ff",
   743 => x"0bd40cd4",
   744 => x"087081ff",
   745 => x"06ff1454",
   746 => x"515171e5",
   747 => x"3870b1d8",
   748 => x"0c028c05",
   749 => x"0d0402fc",
   750 => x"050d81c7",
   751 => x"5181ff0b",
   752 => x"d40cff11",
   753 => x"51708025",
   754 => x"f4380284",
   755 => x"050d0402",
   756 => x"f0050d97",
   757 => x"b62d8fcf",
   758 => x"53805287",
   759 => x"fc80f751",
   760 => x"96c52db1",
   761 => x"d80854b1",
   762 => x"d808812e",
   763 => x"098106a3",
   764 => x"3881ff0b",
   765 => x"d40c820a",
   766 => x"52849c80",
   767 => x"e95196c5",
   768 => x"2db1d808",
   769 => x"8b3881ff",
   770 => x"0bd40c73",
   771 => x"53989904",
   772 => x"97b62dff",
   773 => x"135372c1",
   774 => x"3872b1d8",
   775 => x"0c029005",
   776 => x"0d0402f4",
   777 => x"050d81ff",
   778 => x"0bd40c93",
   779 => x"53805287",
   780 => x"fc80c151",
   781 => x"96c52db1",
   782 => x"d8088b38",
   783 => x"81ff0bd4",
   784 => x"0c815398",
   785 => x"cf0497b6",
   786 => x"2dff1353",
   787 => x"72df3872",
   788 => x"b1d80c02",
   789 => x"8c050d04",
   790 => x"02f0050d",
   791 => x"97b62d83",
   792 => x"aa52849c",
   793 => x"80c85196",
   794 => x"c52db1d8",
   795 => x"08812e09",
   796 => x"81069238",
   797 => x"95f72db1",
   798 => x"d80883ff",
   799 => x"ff065372",
   800 => x"83aa2e97",
   801 => x"3898a22d",
   802 => x"99960481",
   803 => x"549a8504",
   804 => x"aeb45185",
   805 => x"fc2d8054",
   806 => x"9a850481",
   807 => x"ff0bd40c",
   808 => x"b15397cf",
   809 => x"2db1d808",
   810 => x"802e80ca",
   811 => x"38805287",
   812 => x"fc80fa51",
   813 => x"96c52db1",
   814 => x"d808b138",
   815 => x"81ff0bd4",
   816 => x"0cd40853",
   817 => x"81ff0bd4",
   818 => x"0c81ff0b",
   819 => x"d40c81ff",
   820 => x"0bd40c81",
   821 => x"ff0bd40c",
   822 => x"72862a70",
   823 => x"8106b1d8",
   824 => x"08565153",
   825 => x"72802e9d",
   826 => x"38998b04",
   827 => x"b1d80852",
   828 => x"aed0519e",
   829 => x"cb2d7282",
   830 => x"2eff9538",
   831 => x"ff135372",
   832 => x"ffa03872",
   833 => x"5473b1d8",
   834 => x"0c029005",
   835 => x"0d0402f4",
   836 => x"050d810b",
   837 => x"b6b40cd0",
   838 => x"08708f2a",
   839 => x"70810651",
   840 => x"515372f3",
   841 => x"3872d00c",
   842 => x"97b62dae",
   843 => x"dc5185fc",
   844 => x"2dd00870",
   845 => x"8f2a7081",
   846 => x"06515153",
   847 => x"72f33881",
   848 => x"0bd00c80",
   849 => x"e3538052",
   850 => x"84d480c0",
   851 => x"5196c52d",
   852 => x"b1d80881",
   853 => x"2e9a3872",
   854 => x"822e0981",
   855 => x"068c38ae",
   856 => x"f85185fc",
   857 => x"2d80539b",
   858 => x"a504ff13",
   859 => x"5372d738",
   860 => x"98d82db1",
   861 => x"d808b6b4",
   862 => x"0cb1d808",
   863 => x"8b388152",
   864 => x"87fc80d0",
   865 => x"5196c52d",
   866 => x"81ff0bd4",
   867 => x"0cd00870",
   868 => x"8f2a7081",
   869 => x"06515153",
   870 => x"72f33872",
   871 => x"d00c81ff",
   872 => x"0bd40c81",
   873 => x"5372b1d8",
   874 => x"0c028c05",
   875 => x"0d0402e0",
   876 => x"050d797b",
   877 => x"57578058",
   878 => x"81ff0bd4",
   879 => x"0cd00870",
   880 => x"8f2a7081",
   881 => x"06515154",
   882 => x"73f33882",
   883 => x"810bd00c",
   884 => x"81ff0bd4",
   885 => x"0c765287",
   886 => x"fc80d151",
   887 => x"96c52d80",
   888 => x"dbc6df55",
   889 => x"b1d80880",
   890 => x"2e9038b1",
   891 => x"d8085376",
   892 => x"52af9051",
   893 => x"9ecb2d9c",
   894 => x"c80481ff",
   895 => x"0bd40cd4",
   896 => x"087081ff",
   897 => x"06515473",
   898 => x"81fe2e09",
   899 => x"81069d38",
   900 => x"80ff5495",
   901 => x"f72db1d8",
   902 => x"08767084",
   903 => x"05580cff",
   904 => x"14547380",
   905 => x"25ed3881",
   906 => x"589cb204",
   907 => x"ff155574",
   908 => x"c93881ff",
   909 => x"0bd40cd0",
   910 => x"08708f2a",
   911 => x"70810651",
   912 => x"515473f3",
   913 => x"3873d00c",
   914 => x"77b1d80c",
   915 => x"02a0050d",
   916 => x"04b6b408",
   917 => x"b1d80c04",
   918 => x"02e8050d",
   919 => x"80785755",
   920 => x"75708405",
   921 => x"57085380",
   922 => x"5472982a",
   923 => x"73882b54",
   924 => x"5271802e",
   925 => x"a238c008",
   926 => x"70882a70",
   927 => x"81065151",
   928 => x"5170802e",
   929 => x"f13871c0",
   930 => x"0c811581",
   931 => x"15555583",
   932 => x"7425d638",
   933 => x"71ca3874",
   934 => x"b1d80c02",
   935 => x"98050d04",
   936 => x"02f4050d",
   937 => x"7470882a",
   938 => x"83fe8006",
   939 => x"7072982a",
   940 => x"0772882b",
   941 => x"87fc8080",
   942 => x"0673982b",
   943 => x"81f00a06",
   944 => x"71730707",
   945 => x"b1d80c56",
   946 => x"51535102",
   947 => x"8c050d04",
   948 => x"02f8050d",
   949 => x"028e0580",
   950 => x"f52d7488",
   951 => x"2b077083",
   952 => x"ffff06b1",
   953 => x"d80c5102",
   954 => x"88050d04",
   955 => x"02ec050d",
   956 => x"76538055",
   957 => x"7275258b",
   958 => x"38ad5182",
   959 => x"ee2d7209",
   960 => x"81055372",
   961 => x"802eb538",
   962 => x"8754729c",
   963 => x"2a73842b",
   964 => x"54527180",
   965 => x"2e833881",
   966 => x"55897225",
   967 => x"8738b712",
   968 => x"529ea704",
   969 => x"b0125274",
   970 => x"802e8638",
   971 => x"715182ee",
   972 => x"2dff1454",
   973 => x"738025d2",
   974 => x"389ec104",
   975 => x"b05182ee",
   976 => x"2d800bb1",
   977 => x"d80c0294",
   978 => x"050d0402",
   979 => x"c0050d02",
   980 => x"80c40557",
   981 => x"80707870",
   982 => x"84055a08",
   983 => x"72415f5d",
   984 => x"587c7084",
   985 => x"055e085a",
   986 => x"805b7998",
   987 => x"2a7a882b",
   988 => x"5b567586",
   989 => x"38775fa0",
   990 => x"c3047d80",
   991 => x"2e81a238",
   992 => x"805e7580",
   993 => x"e42e8a38",
   994 => x"7580f82e",
   995 => x"09810689",
   996 => x"38768418",
   997 => x"71085e58",
   998 => x"547580e4",
   999 => x"2e9f3875",
  1000 => x"80e4268a",
  1001 => x"387580e3",
  1002 => x"2ebe389f",
  1003 => x"f3047580",
  1004 => x"f32ea338",
  1005 => x"7580f82e",
  1006 => x"89389ff3",
  1007 => x"048a539f",
  1008 => x"c4049053",
  1009 => x"b6b8527b",
  1010 => x"519dec2d",
  1011 => x"b1d808b6",
  1012 => x"b85a55a0",
  1013 => x"83047684",
  1014 => x"18710870",
  1015 => x"545b5854",
  1016 => x"9cd82d80",
  1017 => x"55a08304",
  1018 => x"76841871",
  1019 => x"08585854",
  1020 => x"a0ae04a5",
  1021 => x"5182ee2d",
  1022 => x"755182ee",
  1023 => x"2d821858",
  1024 => x"a0b60474",
  1025 => x"ff165654",
  1026 => x"807425aa",
  1027 => x"38787081",
  1028 => x"055a80f5",
  1029 => x"2d705256",
  1030 => x"82ee2d81",
  1031 => x"1858a083",
  1032 => x"0475a52e",
  1033 => x"09810686",
  1034 => x"38815ea0",
  1035 => x"b6047551",
  1036 => x"82ee2d81",
  1037 => x"1858811b",
  1038 => x"5b837b25",
  1039 => x"feac3875",
  1040 => x"fe9f387e",
  1041 => x"b1d80c02",
  1042 => x"80c0050d",
  1043 => x"0402fc05",
  1044 => x"0d725180",
  1045 => x"710c800b",
  1046 => x"84120c02",
  1047 => x"84050d04",
  1048 => x"02f0050d",
  1049 => x"75700884",
  1050 => x"12085353",
  1051 => x"53ff5471",
  1052 => x"712e9b38",
  1053 => x"84130870",
  1054 => x"8429148b",
  1055 => x"1180f52d",
  1056 => x"84160881",
  1057 => x"11870684",
  1058 => x"180c5256",
  1059 => x"515173b1",
  1060 => x"d80c0290",
  1061 => x"050d0402",
  1062 => x"f8050da4",
  1063 => x"8e2de008",
  1064 => x"708b2a70",
  1065 => x"81065152",
  1066 => x"5270802e",
  1067 => x"9d38b6f8",
  1068 => x"08708429",
  1069 => x"b7800573",
  1070 => x"81ff0671",
  1071 => x"0c5151b6",
  1072 => x"f8088111",
  1073 => x"8706b6f8",
  1074 => x"0c51800b",
  1075 => x"b7a00ca4",
  1076 => x"812da488",
  1077 => x"2d028805",
  1078 => x"0d0402fc",
  1079 => x"050da48e",
  1080 => x"2d810bb7",
  1081 => x"a00ca488",
  1082 => x"2db7a008",
  1083 => x"5170fa38",
  1084 => x"0284050d",
  1085 => x"0402fc05",
  1086 => x"0db6f851",
  1087 => x"a0cd2da1",
  1088 => x"9751a3fd",
  1089 => x"2da3a72d",
  1090 => x"0284050d",
  1091 => x"0402f405",
  1092 => x"0da38f04",
  1093 => x"b1d80881",
  1094 => x"f02e0981",
  1095 => x"06893881",
  1096 => x"0bb1cc0c",
  1097 => x"a38f04b1",
  1098 => x"d80881e0",
  1099 => x"2e098106",
  1100 => x"8938810b",
  1101 => x"b1d00ca3",
  1102 => x"8f04b1d8",
  1103 => x"0852b1d0",
  1104 => x"08802e88",
  1105 => x"38b1d808",
  1106 => x"81800552",
  1107 => x"71842c72",
  1108 => x"8f065353",
  1109 => x"b1cc0880",
  1110 => x"2e993872",
  1111 => x"8429b18c",
  1112 => x"05721381",
  1113 => x"712b7009",
  1114 => x"73080673",
  1115 => x"0c515353",
  1116 => x"a3850472",
  1117 => x"8429b18c",
  1118 => x"05721383",
  1119 => x"712b7208",
  1120 => x"07720c53",
  1121 => x"53800bb1",
  1122 => x"d00c800b",
  1123 => x"b1cc0cb6",
  1124 => x"f851a0e0",
  1125 => x"2db1d808",
  1126 => x"ff24fef8",
  1127 => x"38800bb1",
  1128 => x"d80c028c",
  1129 => x"050d0402",
  1130 => x"f8050db1",
  1131 => x"8c528f51",
  1132 => x"80727084",
  1133 => x"05540cff",
  1134 => x"11517080",
  1135 => x"25f23802",
  1136 => x"88050d04",
  1137 => x"02f0050d",
  1138 => x"7551a48e",
  1139 => x"2d70822c",
  1140 => x"fc06b18c",
  1141 => x"1172109e",
  1142 => x"06710870",
  1143 => x"722a7083",
  1144 => x"0682742b",
  1145 => x"70097406",
  1146 => x"760c5451",
  1147 => x"56575351",
  1148 => x"53a4882d",
  1149 => x"71b1d80c",
  1150 => x"0290050d",
  1151 => x"0471980c",
  1152 => x"04ffb008",
  1153 => x"b1d80c04",
  1154 => x"810bffb0",
  1155 => x"0c04800b",
  1156 => x"ffb00c04",
  1157 => x"02fc050d",
  1158 => x"800bb1d4",
  1159 => x"0c805184",
  1160 => x"e52d0284",
  1161 => x"050d0402",
  1162 => x"f0050db7",
  1163 => x"a8085481",
  1164 => x"f72d800b",
  1165 => x"b7ac0c73",
  1166 => x"08802e80",
  1167 => x"eb38820b",
  1168 => x"b1ec0cb7",
  1169 => x"ac088f06",
  1170 => x"b1e80c73",
  1171 => x"08527181",
  1172 => x"2ea43871",
  1173 => x"832e0981",
  1174 => x"06b93888",
  1175 => x"1480f52d",
  1176 => x"841508af",
  1177 => x"b0535452",
  1178 => x"85fc2d71",
  1179 => x"84291370",
  1180 => x"085252a5",
  1181 => x"9704b7a4",
  1182 => x"08881508",
  1183 => x"2c708106",
  1184 => x"51527180",
  1185 => x"2e8738af",
  1186 => x"b451a590",
  1187 => x"04afb851",
  1188 => x"85fc2d84",
  1189 => x"14085185",
  1190 => x"fc2db7ac",
  1191 => x"088105b7",
  1192 => x"ac0c8c14",
  1193 => x"54a4b704",
  1194 => x"0290050d",
  1195 => x"0471b7a8",
  1196 => x"0ca4a72d",
  1197 => x"b7ac08ff",
  1198 => x"05b7b00c",
  1199 => x"0402f005",
  1200 => x"0d8751a3",
  1201 => x"c42db1d8",
  1202 => x"08812a70",
  1203 => x"81065152",
  1204 => x"71802ea0",
  1205 => x"38a5db04",
  1206 => x"a28d2d87",
  1207 => x"51a3c42d",
  1208 => x"b1d808f4",
  1209 => x"38b1d408",
  1210 => x"813270b1",
  1211 => x"d40c7052",
  1212 => x"5284e52d",
  1213 => x"b1d40896",
  1214 => x"3880da51",
  1215 => x"a3c42d81",
  1216 => x"f551a3c4",
  1217 => x"2d81f251",
  1218 => x"a3c42da8",
  1219 => x"ab0481f5",
  1220 => x"51a3c42d",
  1221 => x"b1d80881",
  1222 => x"2a708106",
  1223 => x"51527180",
  1224 => x"2e8f38b7",
  1225 => x"b0085271",
  1226 => x"802e8638",
  1227 => x"ff12b7b0",
  1228 => x"0c81f251",
  1229 => x"a3c42db1",
  1230 => x"d808812a",
  1231 => x"70810651",
  1232 => x"5271802e",
  1233 => x"9538b7ac",
  1234 => x"08ff05b7",
  1235 => x"b0085452",
  1236 => x"72722586",
  1237 => x"388113b7",
  1238 => x"b00c80da",
  1239 => x"51a3c42d",
  1240 => x"b1d80881",
  1241 => x"2a708106",
  1242 => x"51527180",
  1243 => x"2e80fb38",
  1244 => x"b7a808b7",
  1245 => x"b0085553",
  1246 => x"73802e8a",
  1247 => x"388c13ff",
  1248 => x"155553a6",
  1249 => x"f8047208",
  1250 => x"5271822e",
  1251 => x"a6387182",
  1252 => x"26893871",
  1253 => x"812ea538",
  1254 => x"a7ea0471",
  1255 => x"832ead38",
  1256 => x"71842e09",
  1257 => x"810680c2",
  1258 => x"38881308",
  1259 => x"51a5ad2d",
  1260 => x"a7ea0488",
  1261 => x"13085271",
  1262 => x"2da7ea04",
  1263 => x"810b8814",
  1264 => x"082bb7a4",
  1265 => x"0832b7a4",
  1266 => x"0ca7e704",
  1267 => x"881380f5",
  1268 => x"2d81058b",
  1269 => x"1480f52d",
  1270 => x"53547174",
  1271 => x"24833880",
  1272 => x"54738814",
  1273 => x"81b72da4",
  1274 => x"a72d8054",
  1275 => x"800bb1ec",
  1276 => x"0c738f06",
  1277 => x"b1e80ca0",
  1278 => x"5273b7b0",
  1279 => x"082e0981",
  1280 => x"069838b7",
  1281 => x"ac08ff05",
  1282 => x"74327009",
  1283 => x"81057072",
  1284 => x"079f2a91",
  1285 => x"71315151",
  1286 => x"53537151",
  1287 => x"82ee2d81",
  1288 => x"14548e74",
  1289 => x"25c638b1",
  1290 => x"d4085271",
  1291 => x"b1d80c02",
  1292 => x"90050d04",
  1293 => x"00ffffff",
  1294 => x"ff00ffff",
  1295 => x"ffff00ff",
  1296 => x"ffffff00",
  1297 => x"44495020",
  1298 => x"53776974",
  1299 => x"63686573",
  1300 => x"20100000",
  1301 => x"52657365",
  1302 => x"74000000",
  1303 => x"45786974",
  1304 => x"00000000",
  1305 => x"53442043",
  1306 => x"61726400",
  1307 => x"4a617061",
  1308 => x"6e657365",
  1309 => x"206b6579",
  1310 => x"626f6172",
  1311 => x"64206c61",
  1312 => x"796f7574",
  1313 => x"00000000",
  1314 => x"54757262",
  1315 => x"6f202831",
  1316 => x"302e3734",
  1317 => x"4d487a29",
  1318 => x"00000000",
  1319 => x"4261636b",
  1320 => x"00000000",
  1321 => x"32303438",
  1322 => x"4c422052",
  1323 => x"414d0000",
  1324 => x"34303936",
  1325 => x"4b422052",
  1326 => x"414d0000",
  1327 => x"536c323a",
  1328 => x"204e6f6e",
  1329 => x"65000000",
  1330 => x"536c323a",
  1331 => x"20455345",
  1332 => x"2d534343",
  1333 => x"20314d42",
  1334 => x"2f534343",
  1335 => x"2d490000",
  1336 => x"536c323a",
  1337 => x"20455345",
  1338 => x"2d52414d",
  1339 => x"20314d42",
  1340 => x"2f415343",
  1341 => x"49493800",
  1342 => x"536c323a",
  1343 => x"20455345",
  1344 => x"2d52414d",
  1345 => x"20314d42",
  1346 => x"2f415343",
  1347 => x"49493136",
  1348 => x"00000000",
  1349 => x"536c313a",
  1350 => x"204e6f6e",
  1351 => x"65000000",
  1352 => x"536c313a",
  1353 => x"20455345",
  1354 => x"2d534343",
  1355 => x"20314d42",
  1356 => x"2f534343",
  1357 => x"2d490000",
  1358 => x"536c313a",
  1359 => x"204d6567",
  1360 => x"6152414d",
  1361 => x"00000000",
  1362 => x"56474120",
  1363 => x"2d203331",
  1364 => x"4b487a2c",
  1365 => x"20363048",
  1366 => x"7a000000",
  1367 => x"56474120",
  1368 => x"2d203331",
  1369 => x"4b487a2c",
  1370 => x"20353048",
  1371 => x"7a000000",
  1372 => x"5456202d",
  1373 => x"20343830",
  1374 => x"692c2036",
  1375 => x"30487a00",
  1376 => x"496e6974",
  1377 => x"69616c69",
  1378 => x"7a696e67",
  1379 => x"20534420",
  1380 => x"63617264",
  1381 => x"0a000000",
  1382 => x"53444843",
  1383 => x"20636172",
  1384 => x"64206465",
  1385 => x"74656374",
  1386 => x"65642062",
  1387 => x"7574206e",
  1388 => x"6f740a73",
  1389 => x"7570706f",
  1390 => x"72746564",
  1391 => x"3b206469",
  1392 => x"7361626c",
  1393 => x"696e6720",
  1394 => x"53442063",
  1395 => x"6172640a",
  1396 => x"10204f4b",
  1397 => x"0a000000",
  1398 => x"46617433",
  1399 => x"32206669",
  1400 => x"6c657379",
  1401 => x"7374656d",
  1402 => x"20646574",
  1403 => x"65637465",
  1404 => x"64206275",
  1405 => x"740a6e6f",
  1406 => x"74207375",
  1407 => x"70706f72",
  1408 => x"7465643b",
  1409 => x"20646973",
  1410 => x"61626c69",
  1411 => x"6e672053",
  1412 => x"44206361",
  1413 => x"72640a10",
  1414 => x"204f4b0a",
  1415 => x"00000000",
  1416 => x"54727969",
  1417 => x"6e67204d",
  1418 => x"53583342",
  1419 => x"494f532e",
  1420 => x"5359532e",
  1421 => x"2e2e0a00",
  1422 => x"4d535833",
  1423 => x"42494f53",
  1424 => x"53595300",
  1425 => x"54727969",
  1426 => x"6e672042",
  1427 => x"494f535f",
  1428 => x"4d32502e",
  1429 => x"524f4d2e",
  1430 => x"2e2e0a00",
  1431 => x"42494f53",
  1432 => x"5f4d3250",
  1433 => x"524f4d00",
  1434 => x"4f70656e",
  1435 => x"65642042",
  1436 => x"494f532c",
  1437 => x"206c6f61",
  1438 => x"64696e67",
  1439 => x"2e2e2e0a",
  1440 => x"00000000",
  1441 => x"52656164",
  1442 => x"20626c6f",
  1443 => x"636b2066",
  1444 => x"61696c65",
  1445 => x"640a0000",
  1446 => x"4c6f6164",
  1447 => x"696e6720",
  1448 => x"42494f53",
  1449 => x"20666169",
  1450 => x"6c65640a",
  1451 => x"00000000",
  1452 => x"52656164",
  1453 => x"206f6620",
  1454 => x"4d425220",
  1455 => x"6661696c",
  1456 => x"65640a00",
  1457 => x"46415431",
  1458 => x"36202020",
  1459 => x"00000000",
  1460 => x"46415433",
  1461 => x"32202020",
  1462 => x"00000000",
  1463 => x"25642070",
  1464 => x"61727469",
  1465 => x"74696f6e",
  1466 => x"7320666f",
  1467 => x"756e640a",
  1468 => x"00000000",
  1469 => x"4e6f2070",
  1470 => x"61727469",
  1471 => x"74696f6e",
  1472 => x"20736967",
  1473 => x"6e617475",
  1474 => x"72652066",
  1475 => x"6f756e64",
  1476 => x"0a000000",
  1477 => x"556e7375",
  1478 => x"70706f72",
  1479 => x"74656420",
  1480 => x"70617274",
  1481 => x"6974696f",
  1482 => x"6e207479",
  1483 => x"7065210a",
  1484 => x"00000000",
  1485 => x"53444843",
  1486 => x"20496e69",
  1487 => x"7469616c",
  1488 => x"697a6174",
  1489 => x"696f6e20",
  1490 => x"6572726f",
  1491 => x"72210a00",
  1492 => x"434d4435",
  1493 => x"38202564",
  1494 => x"0a202000",
  1495 => x"496e6974",
  1496 => x"69616c69",
  1497 => x"73696e67",
  1498 => x"20534420",
  1499 => x"63617264",
  1500 => x"2e2e2e0a",
  1501 => x"00000000",
  1502 => x"53442063",
  1503 => x"61726420",
  1504 => x"72657365",
  1505 => x"74206661",
  1506 => x"696c6564",
  1507 => x"210a0000",
  1508 => x"52656164",
  1509 => x"20636f6d",
  1510 => x"6d616e64",
  1511 => x"20666169",
  1512 => x"6c656420",
  1513 => x"61742025",
  1514 => x"64202825",
  1515 => x"64290a00",
  1516 => x"16200000",
  1517 => x"14200000",
  1518 => x"15200000",
  1519 => x"00000002",
  1520 => x"00000004",
  1521 => x"00001444",
  1522 => x"000017f0",
  1523 => x"00000002",
  1524 => x"00001454",
  1525 => x"00000547",
  1526 => x"00000002",
  1527 => x"0000145c",
  1528 => x"00001214",
  1529 => x"00000000",
  1530 => x"00000000",
  1531 => x"00000000",
  1532 => x"00000003",
  1533 => x"00001880",
  1534 => x"00000003",
  1535 => x"00000001",
  1536 => x"00001464",
  1537 => x"00000002",
  1538 => x"00000003",
  1539 => x"00001874",
  1540 => x"00000003",
  1541 => x"00000003",
  1542 => x"00001864",
  1543 => x"00000004",
  1544 => x"00000001",
  1545 => x"0000146c",
  1546 => x"00000006",
  1547 => x"00000001",
  1548 => x"00001488",
  1549 => x"00000007",
  1550 => x"00000003",
  1551 => x"0000185c",
  1552 => x"00000002",
  1553 => x"00000004",
  1554 => x"0000149c",
  1555 => x"000017c0",
  1556 => x"00000000",
  1557 => x"00000000",
  1558 => x"00000000",
  1559 => x"000014a4",
  1560 => x"000014b0",
  1561 => x"000014bc",
  1562 => x"000014c8",
  1563 => x"000014e0",
  1564 => x"000014f8",
  1565 => x"00001514",
  1566 => x"00001520",
  1567 => x"00001538",
  1568 => x"00001548",
  1569 => x"0000155c",
  1570 => x"00001570",
  1571 => x"00000000",
  1572 => x"00000000",
  1573 => x"00000000",
  1574 => x"00000000",
  1575 => x"00000000",
  1576 => x"00000000",
  1577 => x"00000000",
  1578 => x"00000000",
  1579 => x"00000000",
  1580 => x"00000000",
  1581 => x"00000000",
  1582 => x"00000000",
  1583 => x"00000000",
  1584 => x"00000000",
  1585 => x"00000000",
  1586 => x"00000000",
  1587 => x"00000000",
  1588 => x"00000000",
  1589 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

