library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity CharROM_ROM is
generic
	(
		addrbits : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clock : in std_logic;
	address : in std_logic_vector(addrbits-1 downto 0);
	q : out std_logic
);
end CharROM_ROM;

architecture arch of CharROM_ROM is

type rom_type is array(natural range 0 to (2**(addrbits)-1)) of std_logic;

shared variable rom : rom_type :=
(
     0 => '1',
     1 => '0',
     2 => '0',
     3 => '0',
     4 => '0',
     5 => '0',
     6 => '0',
     7 => '0',
     8 => '1',
     9 => '0',
    10 => '0',
    11 => '0',
    12 => '0',
    13 => '0',
    14 => '0',
    15 => '0',
    16 => '1',
    17 => '0',
    18 => '0',
    19 => '0',
    20 => '0',
    21 => '0',
    22 => '0',
    23 => '0',
    24 => '1',
    25 => '0',
    26 => '0',
    27 => '0',
    28 => '0',
    29 => '0',
    30 => '0',
    31 => '0',
    32 => '1',
    33 => '0',
    34 => '0',
    35 => '0',
    36 => '0',
    37 => '0',
    38 => '0',
    39 => '0',
    40 => '1',
    41 => '0',
    42 => '0',
    43 => '0',
    44 => '0',
    45 => '0',
    46 => '0',
    47 => '0',
    48 => '1',
    49 => '0',
    50 => '0',
    51 => '0',
    52 => '0',
    53 => '0',
    54 => '0',
    55 => '0',
    56 => '1',
    57 => '0',
    58 => '0',
    59 => '0',
    60 => '0',
    61 => '0',
    62 => '0',
    63 => '0',
    64 => '1',
    65 => '1',
    66 => '0',
    67 => '0',
    68 => '0',
    69 => '0',
    70 => '0',
    71 => '0',
    72 => '1',
    73 => '1',
    74 => '0',
    75 => '0',
    76 => '0',
    77 => '0',
    78 => '0',
    79 => '0',
    80 => '1',
    81 => '1',
    82 => '0',
    83 => '0',
    84 => '0',
    85 => '0',
    86 => '0',
    87 => '0',
    88 => '1',
    89 => '1',
    90 => '0',
    91 => '0',
    92 => '0',
    93 => '0',
    94 => '0',
    95 => '0',
    96 => '1',
    97 => '1',
    98 => '0',
    99 => '0',
   100 => '0',
   101 => '0',
   102 => '0',
   103 => '0',
   104 => '1',
   105 => '1',
   106 => '0',
   107 => '0',
   108 => '0',
   109 => '0',
   110 => '0',
   111 => '0',
   112 => '1',
   113 => '1',
   114 => '0',
   115 => '0',
   116 => '0',
   117 => '0',
   118 => '0',
   119 => '0',
   120 => '1',
   121 => '1',
   122 => '0',
   123 => '0',
   124 => '0',
   125 => '0',
   126 => '0',
   127 => '0',
   128 => '1',
   129 => '1',
   130 => '1',
   131 => '0',
   132 => '0',
   133 => '0',
   134 => '0',
   135 => '0',
   136 => '1',
   137 => '1',
   138 => '1',
   139 => '0',
   140 => '0',
   141 => '0',
   142 => '0',
   143 => '0',
   144 => '1',
   145 => '1',
   146 => '1',
   147 => '0',
   148 => '0',
   149 => '0',
   150 => '0',
   151 => '0',
   152 => '1',
   153 => '1',
   154 => '1',
   155 => '0',
   156 => '0',
   157 => '0',
   158 => '0',
   159 => '0',
   160 => '1',
   161 => '1',
   162 => '1',
   163 => '0',
   164 => '0',
   165 => '0',
   166 => '0',
   167 => '0',
   168 => '1',
   169 => '1',
   170 => '1',
   171 => '0',
   172 => '0',
   173 => '0',
   174 => '0',
   175 => '0',
   176 => '1',
   177 => '1',
   178 => '1',
   179 => '0',
   180 => '0',
   181 => '0',
   182 => '0',
   183 => '0',
   184 => '1',
   185 => '1',
   186 => '1',
   187 => '0',
   188 => '0',
   189 => '0',
   190 => '0',
   191 => '0',
   192 => '1',
   193 => '1',
   194 => '1',
   195 => '1',
   196 => '0',
   197 => '0',
   198 => '0',
   199 => '0',
   200 => '1',
   201 => '1',
   202 => '1',
   203 => '1',
   204 => '0',
   205 => '0',
   206 => '0',
   207 => '0',
   208 => '1',
   209 => '1',
   210 => '1',
   211 => '1',
   212 => '0',
   213 => '0',
   214 => '0',
   215 => '0',
   216 => '1',
   217 => '1',
   218 => '1',
   219 => '1',
   220 => '0',
   221 => '0',
   222 => '0',
   223 => '0',
   224 => '1',
   225 => '1',
   226 => '1',
   227 => '1',
   228 => '0',
   229 => '0',
   230 => '0',
   231 => '0',
   232 => '1',
   233 => '1',
   234 => '1',
   235 => '1',
   236 => '0',
   237 => '0',
   238 => '0',
   239 => '0',
   240 => '1',
   241 => '1',
   242 => '1',
   243 => '1',
   244 => '0',
   245 => '0',
   246 => '0',
   247 => '0',
   248 => '1',
   249 => '1',
   250 => '1',
   251 => '1',
   252 => '0',
   253 => '0',
   254 => '0',
   255 => '0',
   256 => '1',
   257 => '1',
   258 => '1',
   259 => '1',
   260 => '1',
   261 => '0',
   262 => '0',
   263 => '0',
   264 => '1',
   265 => '1',
   266 => '1',
   267 => '1',
   268 => '1',
   269 => '0',
   270 => '0',
   271 => '0',
   272 => '1',
   273 => '1',
   274 => '1',
   275 => '1',
   276 => '1',
   277 => '0',
   278 => '0',
   279 => '0',
   280 => '1',
   281 => '1',
   282 => '1',
   283 => '1',
   284 => '1',
   285 => '0',
   286 => '0',
   287 => '0',
   288 => '1',
   289 => '1',
   290 => '1',
   291 => '1',
   292 => '1',
   293 => '0',
   294 => '0',
   295 => '0',
   296 => '1',
   297 => '1',
   298 => '1',
   299 => '1',
   300 => '1',
   301 => '0',
   302 => '0',
   303 => '0',
   304 => '1',
   305 => '1',
   306 => '1',
   307 => '1',
   308 => '1',
   309 => '0',
   310 => '0',
   311 => '0',
   312 => '1',
   313 => '1',
   314 => '1',
   315 => '1',
   316 => '1',
   317 => '0',
   318 => '0',
   319 => '0',
   320 => '1',
   321 => '1',
   322 => '1',
   323 => '1',
   324 => '1',
   325 => '1',
   326 => '0',
   327 => '0',
   328 => '1',
   329 => '1',
   330 => '1',
   331 => '1',
   332 => '1',
   333 => '1',
   334 => '0',
   335 => '0',
   336 => '1',
   337 => '1',
   338 => '1',
   339 => '1',
   340 => '1',
   341 => '1',
   342 => '0',
   343 => '0',
   344 => '1',
   345 => '1',
   346 => '1',
   347 => '1',
   348 => '1',
   349 => '1',
   350 => '0',
   351 => '0',
   352 => '1',
   353 => '1',
   354 => '1',
   355 => '1',
   356 => '1',
   357 => '1',
   358 => '0',
   359 => '0',
   360 => '1',
   361 => '1',
   362 => '1',
   363 => '1',
   364 => '1',
   365 => '1',
   366 => '0',
   367 => '0',
   368 => '1',
   369 => '1',
   370 => '1',
   371 => '1',
   372 => '1',
   373 => '1',
   374 => '0',
   375 => '0',
   376 => '1',
   377 => '1',
   378 => '1',
   379 => '1',
   380 => '1',
   381 => '1',
   382 => '0',
   383 => '0',
   384 => '1',
   385 => '1',
   386 => '1',
   387 => '1',
   388 => '1',
   389 => '1',
   390 => '1',
   391 => '0',
   392 => '1',
   393 => '1',
   394 => '1',
   395 => '1',
   396 => '1',
   397 => '1',
   398 => '1',
   399 => '0',
   400 => '1',
   401 => '1',
   402 => '1',
   403 => '1',
   404 => '1',
   405 => '1',
   406 => '1',
   407 => '0',
   408 => '1',
   409 => '1',
   410 => '1',
   411 => '1',
   412 => '1',
   413 => '1',
   414 => '1',
   415 => '0',
   416 => '1',
   417 => '1',
   418 => '1',
   419 => '1',
   420 => '1',
   421 => '1',
   422 => '1',
   423 => '0',
   424 => '1',
   425 => '1',
   426 => '1',
   427 => '1',
   428 => '1',
   429 => '1',
   430 => '1',
   431 => '0',
   432 => '1',
   433 => '1',
   434 => '1',
   435 => '1',
   436 => '1',
   437 => '1',
   438 => '1',
   439 => '0',
   440 => '1',
   441 => '1',
   442 => '1',
   443 => '1',
   444 => '1',
   445 => '1',
   446 => '1',
   447 => '0',
   448 => '1',
   449 => '1',
   450 => '1',
   451 => '1',
   452 => '1',
   453 => '1',
   454 => '1',
   455 => '1',
   456 => '1',
   457 => '1',
   458 => '1',
   459 => '1',
   460 => '1',
   461 => '1',
   462 => '1',
   463 => '1',
   464 => '1',
   465 => '1',
   466 => '1',
   467 => '1',
   468 => '1',
   469 => '1',
   470 => '1',
   471 => '1',
   472 => '1',
   473 => '1',
   474 => '1',
   475 => '1',
   476 => '1',
   477 => '1',
   478 => '1',
   479 => '1',
   480 => '1',
   481 => '1',
   482 => '1',
   483 => '1',
   484 => '1',
   485 => '1',
   486 => '1',
   487 => '1',
   488 => '1',
   489 => '1',
   490 => '1',
   491 => '1',
   492 => '1',
   493 => '1',
   494 => '1',
   495 => '1',
   496 => '1',
   497 => '1',
   498 => '1',
   499 => '1',
   500 => '1',
   501 => '1',
   502 => '1',
   503 => '1',
   504 => '1',
   505 => '1',
   506 => '1',
   507 => '1',
   508 => '1',
   509 => '1',
   510 => '1',
   511 => '1',
   512 => '0',
   513 => '0',
   514 => '0',
   515 => '0',
   516 => '0',
   517 => '0',
   518 => '0',
   519 => '1',
   520 => '0',
   521 => '0',
   522 => '0',
   523 => '0',
   524 => '0',
   525 => '0',
   526 => '0',
   527 => '1',
   528 => '0',
   529 => '0',
   530 => '0',
   531 => '0',
   532 => '0',
   533 => '0',
   534 => '0',
   535 => '1',
   536 => '0',
   537 => '0',
   538 => '0',
   539 => '0',
   540 => '0',
   541 => '0',
   542 => '0',
   543 => '1',
   544 => '0',
   545 => '0',
   546 => '0',
   547 => '0',
   548 => '0',
   549 => '0',
   550 => '0',
   551 => '1',
   552 => '0',
   553 => '0',
   554 => '0',
   555 => '0',
   556 => '0',
   557 => '0',
   558 => '0',
   559 => '1',
   560 => '0',
   561 => '0',
   562 => '0',
   563 => '0',
   564 => '0',
   565 => '0',
   566 => '0',
   567 => '1',
   568 => '0',
   569 => '0',
   570 => '0',
   571 => '0',
   572 => '0',
   573 => '0',
   574 => '0',
   575 => '1',
   576 => '0',
   577 => '0',
   578 => '0',
   579 => '0',
   580 => '0',
   581 => '0',
   582 => '1',
   583 => '1',
   584 => '0',
   585 => '0',
   586 => '0',
   587 => '0',
   588 => '0',
   589 => '0',
   590 => '1',
   591 => '1',
   592 => '0',
   593 => '0',
   594 => '0',
   595 => '0',
   596 => '0',
   597 => '0',
   598 => '1',
   599 => '1',
   600 => '0',
   601 => '0',
   602 => '0',
   603 => '0',
   604 => '0',
   605 => '0',
   606 => '1',
   607 => '1',
   608 => '0',
   609 => '0',
   610 => '0',
   611 => '0',
   612 => '0',
   613 => '0',
   614 => '1',
   615 => '1',
   616 => '0',
   617 => '0',
   618 => '0',
   619 => '0',
   620 => '0',
   621 => '0',
   622 => '1',
   623 => '1',
   624 => '0',
   625 => '0',
   626 => '0',
   627 => '0',
   628 => '0',
   629 => '0',
   630 => '1',
   631 => '1',
   632 => '0',
   633 => '0',
   634 => '0',
   635 => '0',
   636 => '0',
   637 => '0',
   638 => '1',
   639 => '1',
   640 => '0',
   641 => '0',
   642 => '0',
   643 => '0',
   644 => '0',
   645 => '1',
   646 => '1',
   647 => '1',
   648 => '0',
   649 => '0',
   650 => '0',
   651 => '0',
   652 => '0',
   653 => '1',
   654 => '1',
   655 => '1',
   656 => '0',
   657 => '0',
   658 => '0',
   659 => '0',
   660 => '0',
   661 => '1',
   662 => '1',
   663 => '1',
   664 => '0',
   665 => '0',
   666 => '0',
   667 => '0',
   668 => '0',
   669 => '1',
   670 => '1',
   671 => '1',
   672 => '0',
   673 => '0',
   674 => '0',
   675 => '0',
   676 => '0',
   677 => '1',
   678 => '1',
   679 => '1',
   680 => '0',
   681 => '0',
   682 => '0',
   683 => '0',
   684 => '0',
   685 => '1',
   686 => '1',
   687 => '1',
   688 => '0',
   689 => '0',
   690 => '0',
   691 => '0',
   692 => '0',
   693 => '1',
   694 => '1',
   695 => '1',
   696 => '0',
   697 => '0',
   698 => '0',
   699 => '0',
   700 => '0',
   701 => '1',
   702 => '1',
   703 => '1',
   704 => '0',
   705 => '0',
   706 => '0',
   707 => '0',
   708 => '1',
   709 => '1',
   710 => '1',
   711 => '1',
   712 => '0',
   713 => '0',
   714 => '0',
   715 => '0',
   716 => '1',
   717 => '1',
   718 => '1',
   719 => '1',
   720 => '0',
   721 => '0',
   722 => '0',
   723 => '0',
   724 => '1',
   725 => '1',
   726 => '1',
   727 => '1',
   728 => '0',
   729 => '0',
   730 => '0',
   731 => '0',
   732 => '1',
   733 => '1',
   734 => '1',
   735 => '1',
   736 => '0',
   737 => '0',
   738 => '0',
   739 => '0',
   740 => '1',
   741 => '1',
   742 => '1',
   743 => '1',
   744 => '0',
   745 => '0',
   746 => '0',
   747 => '0',
   748 => '1',
   749 => '1',
   750 => '1',
   751 => '1',
   752 => '0',
   753 => '0',
   754 => '0',
   755 => '0',
   756 => '1',
   757 => '1',
   758 => '1',
   759 => '1',
   760 => '0',
   761 => '0',
   762 => '0',
   763 => '0',
   764 => '1',
   765 => '1',
   766 => '1',
   767 => '1',
   768 => '0',
   769 => '0',
   770 => '0',
   771 => '1',
   772 => '1',
   773 => '1',
   774 => '1',
   775 => '1',
   776 => '0',
   777 => '0',
   778 => '0',
   779 => '1',
   780 => '1',
   781 => '1',
   782 => '1',
   783 => '1',
   784 => '0',
   785 => '0',
   786 => '0',
   787 => '1',
   788 => '1',
   789 => '1',
   790 => '1',
   791 => '1',
   792 => '0',
   793 => '0',
   794 => '0',
   795 => '1',
   796 => '1',
   797 => '1',
   798 => '1',
   799 => '1',
   800 => '0',
   801 => '0',
   802 => '0',
   803 => '1',
   804 => '1',
   805 => '1',
   806 => '1',
   807 => '1',
   808 => '0',
   809 => '0',
   810 => '0',
   811 => '1',
   812 => '1',
   813 => '1',
   814 => '1',
   815 => '1',
   816 => '0',
   817 => '0',
   818 => '0',
   819 => '1',
   820 => '1',
   821 => '1',
   822 => '1',
   823 => '1',
   824 => '0',
   825 => '0',
   826 => '0',
   827 => '1',
   828 => '1',
   829 => '1',
   830 => '1',
   831 => '1',
   832 => '0',
   833 => '0',
   834 => '1',
   835 => '1',
   836 => '1',
   837 => '1',
   838 => '1',
   839 => '1',
   840 => '0',
   841 => '0',
   842 => '1',
   843 => '1',
   844 => '1',
   845 => '1',
   846 => '1',
   847 => '1',
   848 => '0',
   849 => '0',
   850 => '1',
   851 => '1',
   852 => '1',
   853 => '1',
   854 => '1',
   855 => '1',
   856 => '0',
   857 => '0',
   858 => '1',
   859 => '1',
   860 => '1',
   861 => '1',
   862 => '1',
   863 => '1',
   864 => '0',
   865 => '0',
   866 => '1',
   867 => '1',
   868 => '1',
   869 => '1',
   870 => '1',
   871 => '1',
   872 => '0',
   873 => '0',
   874 => '1',
   875 => '1',
   876 => '1',
   877 => '1',
   878 => '1',
   879 => '1',
   880 => '0',
   881 => '0',
   882 => '1',
   883 => '1',
   884 => '1',
   885 => '1',
   886 => '1',
   887 => '1',
   888 => '0',
   889 => '0',
   890 => '1',
   891 => '1',
   892 => '1',
   893 => '1',
   894 => '1',
   895 => '1',
   896 => '0',
   897 => '1',
   898 => '1',
   899 => '1',
   900 => '1',
   901 => '1',
   902 => '1',
   903 => '1',
   904 => '0',
   905 => '1',
   906 => '1',
   907 => '1',
   908 => '1',
   909 => '1',
   910 => '1',
   911 => '1',
   912 => '0',
   913 => '1',
   914 => '1',
   915 => '1',
   916 => '1',
   917 => '1',
   918 => '1',
   919 => '1',
   920 => '0',
   921 => '1',
   922 => '1',
   923 => '1',
   924 => '1',
   925 => '1',
   926 => '1',
   927 => '1',
   928 => '0',
   929 => '1',
   930 => '1',
   931 => '1',
   932 => '1',
   933 => '1',
   934 => '1',
   935 => '1',
   936 => '0',
   937 => '1',
   938 => '1',
   939 => '1',
   940 => '1',
   941 => '1',
   942 => '1',
   943 => '1',
   944 => '0',
   945 => '1',
   946 => '1',
   947 => '1',
   948 => '1',
   949 => '1',
   950 => '1',
   951 => '1',
   952 => '0',
   953 => '1',
   954 => '1',
   955 => '1',
   956 => '1',
   957 => '1',
   958 => '1',
   959 => '1',
   960 => '1',
   961 => '1',
   962 => '1',
   963 => '1',
   964 => '1',
   965 => '1',
   966 => '1',
   967 => '1',
   968 => '1',
   969 => '1',
   970 => '1',
   971 => '1',
   972 => '1',
   973 => '1',
   974 => '1',
   975 => '1',
   976 => '1',
   977 => '1',
   978 => '1',
   979 => '1',
   980 => '1',
   981 => '1',
   982 => '1',
   983 => '1',
   984 => '1',
   985 => '1',
   986 => '1',
   987 => '1',
   988 => '1',
   989 => '1',
   990 => '1',
   991 => '1',
   992 => '1',
   993 => '1',
   994 => '1',
   995 => '1',
   996 => '1',
   997 => '1',
   998 => '1',
   999 => '1',
  1000 => '1',
  1001 => '1',
  1002 => '1',
  1003 => '1',
  1004 => '1',
  1005 => '1',
  1006 => '1',
  1007 => '1',
  1008 => '1',
  1009 => '1',
  1010 => '1',
  1011 => '1',
  1012 => '1',
  1013 => '1',
  1014 => '1',
  1015 => '1',
  1016 => '1',
  1017 => '1',
  1018 => '1',
  1019 => '1',
  1020 => '1',
  1021 => '1',
  1022 => '1',
  1023 => '1',
  1024 => '0',
  1025 => '0',
  1026 => '0',
  1027 => '0',
  1028 => '0',
  1029 => '0',
  1030 => '0',
  1031 => '0',
  1032 => '0',
  1033 => '1',
  1034 => '0',
  1035 => '0',
  1036 => '0',
  1037 => '0',
  1038 => '0',
  1039 => '0',
  1040 => '0',
  1041 => '1',
  1042 => '1',
  1043 => '1',
  1044 => '0',
  1045 => '0',
  1046 => '0',
  1047 => '0',
  1048 => '0',
  1049 => '1',
  1050 => '1',
  1051 => '1',
  1052 => '1',
  1053 => '1',
  1054 => '0',
  1055 => '0',
  1056 => '0',
  1057 => '1',
  1058 => '1',
  1059 => '1',
  1060 => '1',
  1061 => '1',
  1062 => '0',
  1063 => '0',
  1064 => '0',
  1065 => '1',
  1066 => '1',
  1067 => '1',
  1068 => '0',
  1069 => '0',
  1070 => '0',
  1071 => '0',
  1072 => '0',
  1073 => '1',
  1074 => '0',
  1075 => '0',
  1076 => '0',
  1077 => '0',
  1078 => '0',
  1079 => '0',
  1080 => '0',
  1081 => '0',
  1082 => '0',
  1083 => '0',
  1084 => '0',
  1085 => '0',
  1086 => '0',
  1087 => '0',
  1088 => '0',
  1089 => '0',
  1090 => '0',
  1091 => '0',
  1092 => '0',
  1093 => '0',
  1094 => '0',
  1095 => '0',
  1096 => '0',
  1097 => '0',
  1098 => '0',
  1099 => '0',
  1100 => '0',
  1101 => '0',
  1102 => '1',
  1103 => '0',
  1104 => '0',
  1105 => '0',
  1106 => '0',
  1107 => '0',
  1108 => '1',
  1109 => '1',
  1110 => '1',
  1111 => '0',
  1112 => '0',
  1113 => '0',
  1114 => '1',
  1115 => '1',
  1116 => '1',
  1117 => '1',
  1118 => '1',
  1119 => '0',
  1120 => '0',
  1121 => '0',
  1122 => '1',
  1123 => '1',
  1124 => '1',
  1125 => '1',
  1126 => '1',
  1127 => '0',
  1128 => '0',
  1129 => '0',
  1130 => '0',
  1131 => '0',
  1132 => '1',
  1133 => '1',
  1134 => '1',
  1135 => '0',
  1136 => '0',
  1137 => '0',
  1138 => '0',
  1139 => '0',
  1140 => '0',
  1141 => '0',
  1142 => '1',
  1143 => '0',
  1144 => '0',
  1145 => '0',
  1146 => '0',
  1147 => '0',
  1148 => '0',
  1149 => '0',
  1150 => '0',
  1151 => '0',
  1152 => '0',
  1153 => '0',
  1154 => '0',
  1155 => '0',
  1156 => '0',
  1157 => '0',
  1158 => '0',
  1159 => '0',
  1160 => '0',
  1161 => '0',
  1162 => '0',
  1163 => '1',
  1164 => '1',
  1165 => '0',
  1166 => '0',
  1167 => '0',
  1168 => '0',
  1169 => '0',
  1170 => '0',
  1171 => '1',
  1172 => '1',
  1173 => '0',
  1174 => '0',
  1175 => '0',
  1176 => '0',
  1177 => '0',
  1178 => '1',
  1179 => '1',
  1180 => '1',
  1181 => '1',
  1182 => '0',
  1183 => '0',
  1184 => '0',
  1185 => '0',
  1186 => '1',
  1187 => '1',
  1188 => '1',
  1189 => '1',
  1190 => '0',
  1191 => '0',
  1192 => '0',
  1193 => '1',
  1194 => '1',
  1195 => '1',
  1196 => '1',
  1197 => '1',
  1198 => '1',
  1199 => '0',
  1200 => '0',
  1201 => '1',
  1202 => '1',
  1203 => '1',
  1204 => '1',
  1205 => '1',
  1206 => '1',
  1207 => '0',
  1208 => '0',
  1209 => '0',
  1210 => '0',
  1211 => '0',
  1212 => '0',
  1213 => '0',
  1214 => '0',
  1215 => '0',
  1216 => '0',
  1217 => '0',
  1218 => '0',
  1219 => '0',
  1220 => '0',
  1221 => '0',
  1222 => '0',
  1223 => '0',
  1224 => '0',
  1225 => '1',
  1226 => '1',
  1227 => '1',
  1228 => '1',
  1229 => '1',
  1230 => '1',
  1231 => '0',
  1232 => '0',
  1233 => '1',
  1234 => '1',
  1235 => '1',
  1236 => '1',
  1237 => '1',
  1238 => '1',
  1239 => '0',
  1240 => '0',
  1241 => '0',
  1242 => '1',
  1243 => '1',
  1244 => '1',
  1245 => '1',
  1246 => '0',
  1247 => '0',
  1248 => '0',
  1249 => '0',
  1250 => '1',
  1251 => '1',
  1252 => '1',
  1253 => '1',
  1254 => '0',
  1255 => '0',
  1256 => '0',
  1257 => '0',
  1258 => '0',
  1259 => '1',
  1260 => '1',
  1261 => '0',
  1262 => '0',
  1263 => '0',
  1264 => '0',
  1265 => '0',
  1266 => '0',
  1267 => '1',
  1268 => '1',
  1269 => '0',
  1270 => '0',
  1271 => '0',
  1272 => '0',
  1273 => '0',
  1274 => '0',
  1275 => '0',
  1276 => '0',
  1277 => '0',
  1278 => '0',
  1279 => '0',
  1280 => '0',
  1281 => '0',
  1282 => '0',
  1283 => '0',
  1284 => '0',
  1285 => '0',
  1286 => '0',
  1287 => '0',
  1288 => '0',
  1289 => '0',
  1290 => '0',
  1291 => '0',
  1292 => '0',
  1293 => '1',
  1294 => '1',
  1295 => '0',
  1296 => '0',
  1297 => '0',
  1298 => '0',
  1299 => '0',
  1300 => '0',
  1301 => '1',
  1302 => '1',
  1303 => '0',
  1304 => '0',
  1305 => '0',
  1306 => '0',
  1307 => '0',
  1308 => '1',
  1309 => '1',
  1310 => '0',
  1311 => '0',
  1312 => '1',
  1313 => '1',
  1314 => '0',
  1315 => '0',
  1316 => '1',
  1317 => '1',
  1318 => '0',
  1319 => '0',
  1320 => '0',
  1321 => '1',
  1322 => '1',
  1323 => '1',
  1324 => '1',
  1325 => '0',
  1326 => '0',
  1327 => '0',
  1328 => '0',
  1329 => '0',
  1330 => '1',
  1331 => '1',
  1332 => '1',
  1333 => '0',
  1334 => '0',
  1335 => '0',
  1336 => '0',
  1337 => '0',
  1338 => '0',
  1339 => '0',
  1340 => '0',
  1341 => '0',
  1342 => '0',
  1343 => '0',
  1344 => '0',
  1345 => '0',
  1346 => '0',
  1347 => '0',
  1348 => '0',
  1349 => '0',
  1350 => '0',
  1351 => '0',
  1352 => '1',
  1353 => '1',
  1354 => '0',
  1355 => '0',
  1356 => '0',
  1357 => '1',
  1358 => '1',
  1359 => '0',
  1360 => '0',
  1361 => '1',
  1362 => '1',
  1363 => '0',
  1364 => '1',
  1365 => '1',
  1366 => '0',
  1367 => '0',
  1368 => '0',
  1369 => '0',
  1370 => '1',
  1371 => '1',
  1372 => '1',
  1373 => '0',
  1374 => '0',
  1375 => '0',
  1376 => '0',
  1377 => '0',
  1378 => '1',
  1379 => '1',
  1380 => '1',
  1381 => '0',
  1382 => '0',
  1383 => '0',
  1384 => '0',
  1385 => '1',
  1386 => '1',
  1387 => '0',
  1388 => '1',
  1389 => '1',
  1390 => '0',
  1391 => '0',
  1392 => '1',
  1393 => '1',
  1394 => '0',
  1395 => '0',
  1396 => '0',
  1397 => '1',
  1398 => '1',
  1399 => '0',
  1400 => '0',
  1401 => '0',
  1402 => '0',
  1403 => '0',
  1404 => '0',
  1405 => '0',
  1406 => '0',
  1407 => '0',
  1408 => '0',
  1409 => '0',
  1410 => '0',
  1411 => '1',
  1412 => '1',
  1413 => '0',
  1414 => '0',
  1415 => '0',
  1416 => '1',
  1417 => '0',
  1418 => '1',
  1419 => '1',
  1420 => '1',
  1421 => '1',
  1422 => '0',
  1423 => '0',
  1424 => '1',
  1425 => '1',
  1426 => '1',
  1427 => '0',
  1428 => '0',
  1429 => '1',
  1430 => '1',
  1431 => '0',
  1432 => '1',
  1433 => '1',
  1434 => '0',
  1435 => '0',
  1436 => '0',
  1437 => '0',
  1438 => '1',
  1439 => '0',
  1440 => '1',
  1441 => '1',
  1442 => '1',
  1443 => '0',
  1444 => '0',
  1445 => '1',
  1446 => '1',
  1447 => '0',
  1448 => '0',
  1449 => '0',
  1450 => '0',
  1451 => '0',
  1452 => '1',
  1453 => '1',
  1454 => '0',
  1455 => '0',
  1456 => '0',
  1457 => '0',
  1458 => '1',
  1459 => '1',
  1460 => '1',
  1461 => '0',
  1462 => '0',
  1463 => '0',
  1464 => '0',
  1465 => '0',
  1466 => '0',
  1467 => '0',
  1468 => '0',
  1469 => '0',
  1470 => '0',
  1471 => '0',
  1472 => '0',
  1473 => '0',
  1474 => '0',
  1475 => '0',
  1476 => '0',
  1477 => '0',
  1478 => '0',
  1479 => '0',
  1480 => '0',
  1481 => '0',
  1482 => '0',
  1483 => '0',
  1484 => '0',
  1485 => '0',
  1486 => '0',
  1487 => '0',
  1488 => '0',
  1489 => '0',
  1490 => '0',
  1491 => '0',
  1492 => '0',
  1493 => '0',
  1494 => '0',
  1495 => '0',
  1496 => '0',
  1497 => '0',
  1498 => '0',
  1499 => '0',
  1500 => '0',
  1501 => '0',
  1502 => '0',
  1503 => '0',
  1504 => '0',
  1505 => '0',
  1506 => '0',
  1507 => '0',
  1508 => '0',
  1509 => '0',
  1510 => '0',
  1511 => '0',
  1512 => '0',
  1513 => '0',
  1514 => '0',
  1515 => '0',
  1516 => '0',
  1517 => '0',
  1518 => '0',
  1519 => '0',
  1520 => '0',
  1521 => '0',
  1522 => '0',
  1523 => '0',
  1524 => '0',
  1525 => '0',
  1526 => '0',
  1527 => '0',
  1528 => '0',
  1529 => '0',
  1530 => '0',
  1531 => '0',
  1532 => '0',
  1533 => '0',
  1534 => '0',
  1535 => '0',
  1536 => '0',
  1537 => '0',
  1538 => '0',
  1539 => '0',
  1540 => '0',
  1541 => '0',
  1542 => '0',
  1543 => '0',
  1544 => '0',
  1545 => '0',
  1546 => '0',
  1547 => '0',
  1548 => '0',
  1549 => '0',
  1550 => '0',
  1551 => '0',
  1552 => '0',
  1553 => '0',
  1554 => '0',
  1555 => '0',
  1556 => '0',
  1557 => '0',
  1558 => '0',
  1559 => '0',
  1560 => '0',
  1561 => '0',
  1562 => '0',
  1563 => '0',
  1564 => '0',
  1565 => '0',
  1566 => '0',
  1567 => '0',
  1568 => '0',
  1569 => '0',
  1570 => '0',
  1571 => '0',
  1572 => '0',
  1573 => '0',
  1574 => '0',
  1575 => '0',
  1576 => '0',
  1577 => '0',
  1578 => '0',
  1579 => '0',
  1580 => '0',
  1581 => '0',
  1582 => '0',
  1583 => '0',
  1584 => '0',
  1585 => '0',
  1586 => '0',
  1587 => '0',
  1588 => '0',
  1589 => '0',
  1590 => '0',
  1591 => '0',
  1592 => '0',
  1593 => '0',
  1594 => '0',
  1595 => '0',
  1596 => '0',
  1597 => '0',
  1598 => '0',
  1599 => '0',
  1600 => '0',
  1601 => '0',
  1602 => '0',
  1603 => '0',
  1604 => '0',
  1605 => '0',
  1606 => '0',
  1607 => '0',
  1608 => '0',
  1609 => '0',
  1610 => '0',
  1611 => '0',
  1612 => '0',
  1613 => '0',
  1614 => '0',
  1615 => '0',
  1616 => '0',
  1617 => '0',
  1618 => '0',
  1619 => '0',
  1620 => '0',
  1621 => '0',
  1622 => '0',
  1623 => '0',
  1624 => '0',
  1625 => '0',
  1626 => '0',
  1627 => '0',
  1628 => '0',
  1629 => '0',
  1630 => '0',
  1631 => '0',
  1632 => '0',
  1633 => '0',
  1634 => '0',
  1635 => '0',
  1636 => '0',
  1637 => '0',
  1638 => '0',
  1639 => '0',
  1640 => '0',
  1641 => '0',
  1642 => '0',
  1643 => '0',
  1644 => '0',
  1645 => '0',
  1646 => '0',
  1647 => '0',
  1648 => '0',
  1649 => '0',
  1650 => '0',
  1651 => '0',
  1652 => '0',
  1653 => '0',
  1654 => '0',
  1655 => '0',
  1656 => '0',
  1657 => '0',
  1658 => '0',
  1659 => '0',
  1660 => '0',
  1661 => '0',
  1662 => '0',
  1663 => '0',
  1664 => '0',
  1665 => '0',
  1666 => '0',
  1667 => '0',
  1668 => '0',
  1669 => '0',
  1670 => '0',
  1671 => '0',
  1672 => '0',
  1673 => '0',
  1674 => '0',
  1675 => '0',
  1676 => '0',
  1677 => '0',
  1678 => '0',
  1679 => '0',
  1680 => '0',
  1681 => '0',
  1682 => '0',
  1683 => '0',
  1684 => '0',
  1685 => '0',
  1686 => '0',
  1687 => '0',
  1688 => '0',
  1689 => '0',
  1690 => '0',
  1691 => '0',
  1692 => '0',
  1693 => '0',
  1694 => '0',
  1695 => '0',
  1696 => '0',
  1697 => '0',
  1698 => '0',
  1699 => '0',
  1700 => '0',
  1701 => '0',
  1702 => '0',
  1703 => '0',
  1704 => '0',
  1705 => '0',
  1706 => '0',
  1707 => '0',
  1708 => '0',
  1709 => '0',
  1710 => '0',
  1711 => '0',
  1712 => '0',
  1713 => '0',
  1714 => '0',
  1715 => '0',
  1716 => '0',
  1717 => '0',
  1718 => '0',
  1719 => '0',
  1720 => '0',
  1721 => '0',
  1722 => '0',
  1723 => '0',
  1724 => '0',
  1725 => '0',
  1726 => '0',
  1727 => '0',
  1728 => '0',
  1729 => '0',
  1730 => '0',
  1731 => '0',
  1732 => '0',
  1733 => '0',
  1734 => '0',
  1735 => '0',
  1736 => '0',
  1737 => '0',
  1738 => '0',
  1739 => '0',
  1740 => '0',
  1741 => '0',
  1742 => '0',
  1743 => '0',
  1744 => '0',
  1745 => '0',
  1746 => '0',
  1747 => '0',
  1748 => '0',
  1749 => '0',
  1750 => '0',
  1751 => '0',
  1752 => '0',
  1753 => '0',
  1754 => '0',
  1755 => '0',
  1756 => '0',
  1757 => '0',
  1758 => '0',
  1759 => '0',
  1760 => '0',
  1761 => '0',
  1762 => '0',
  1763 => '0',
  1764 => '0',
  1765 => '0',
  1766 => '0',
  1767 => '0',
  1768 => '0',
  1769 => '0',
  1770 => '0',
  1771 => '0',
  1772 => '0',
  1773 => '0',
  1774 => '0',
  1775 => '0',
  1776 => '0',
  1777 => '0',
  1778 => '0',
  1779 => '0',
  1780 => '0',
  1781 => '0',
  1782 => '0',
  1783 => '0',
  1784 => '0',
  1785 => '0',
  1786 => '0',
  1787 => '0',
  1788 => '0',
  1789 => '0',
  1790 => '0',
  1791 => '0',
  1792 => '0',
  1793 => '0',
  1794 => '0',
  1795 => '0',
  1796 => '0',
  1797 => '0',
  1798 => '0',
  1799 => '0',
  1800 => '0',
  1801 => '0',
  1802 => '0',
  1803 => '0',
  1804 => '0',
  1805 => '0',
  1806 => '0',
  1807 => '0',
  1808 => '0',
  1809 => '0',
  1810 => '0',
  1811 => '0',
  1812 => '0',
  1813 => '0',
  1814 => '0',
  1815 => '0',
  1816 => '0',
  1817 => '0',
  1818 => '0',
  1819 => '0',
  1820 => '0',
  1821 => '0',
  1822 => '0',
  1823 => '0',
  1824 => '0',
  1825 => '0',
  1826 => '0',
  1827 => '0',
  1828 => '0',
  1829 => '0',
  1830 => '0',
  1831 => '0',
  1832 => '0',
  1833 => '0',
  1834 => '0',
  1835 => '0',
  1836 => '0',
  1837 => '0',
  1838 => '0',
  1839 => '0',
  1840 => '0',
  1841 => '0',
  1842 => '0',
  1843 => '0',
  1844 => '0',
  1845 => '0',
  1846 => '0',
  1847 => '0',
  1848 => '0',
  1849 => '0',
  1850 => '0',
  1851 => '0',
  1852 => '0',
  1853 => '0',
  1854 => '0',
  1855 => '0',
  1856 => '0',
  1857 => '0',
  1858 => '0',
  1859 => '0',
  1860 => '0',
  1861 => '0',
  1862 => '0',
  1863 => '0',
  1864 => '0',
  1865 => '0',
  1866 => '0',
  1867 => '0',
  1868 => '0',
  1869 => '0',
  1870 => '0',
  1871 => '0',
  1872 => '0',
  1873 => '0',
  1874 => '0',
  1875 => '0',
  1876 => '0',
  1877 => '0',
  1878 => '0',
  1879 => '0',
  1880 => '0',
  1881 => '0',
  1882 => '0',
  1883 => '0',
  1884 => '0',
  1885 => '0',
  1886 => '0',
  1887 => '0',
  1888 => '0',
  1889 => '0',
  1890 => '0',
  1891 => '0',
  1892 => '0',
  1893 => '0',
  1894 => '0',
  1895 => '0',
  1896 => '0',
  1897 => '0',
  1898 => '0',
  1899 => '0',
  1900 => '0',
  1901 => '0',
  1902 => '0',
  1903 => '0',
  1904 => '0',
  1905 => '0',
  1906 => '0',
  1907 => '0',
  1908 => '0',
  1909 => '0',
  1910 => '0',
  1911 => '0',
  1912 => '0',
  1913 => '0',
  1914 => '0',
  1915 => '0',
  1916 => '0',
  1917 => '0',
  1918 => '0',
  1919 => '0',
  1920 => '0',
  1921 => '0',
  1922 => '0',
  1923 => '0',
  1924 => '0',
  1925 => '0',
  1926 => '0',
  1927 => '0',
  1928 => '0',
  1929 => '0',
  1930 => '0',
  1931 => '0',
  1932 => '0',
  1933 => '0',
  1934 => '0',
  1935 => '0',
  1936 => '0',
  1937 => '0',
  1938 => '0',
  1939 => '0',
  1940 => '0',
  1941 => '0',
  1942 => '0',
  1943 => '0',
  1944 => '0',
  1945 => '0',
  1946 => '0',
  1947 => '0',
  1948 => '0',
  1949 => '0',
  1950 => '0',
  1951 => '0',
  1952 => '0',
  1953 => '0',
  1954 => '0',
  1955 => '0',
  1956 => '0',
  1957 => '0',
  1958 => '0',
  1959 => '0',
  1960 => '0',
  1961 => '0',
  1962 => '0',
  1963 => '0',
  1964 => '0',
  1965 => '0',
  1966 => '0',
  1967 => '0',
  1968 => '0',
  1969 => '0',
  1970 => '0',
  1971 => '0',
  1972 => '0',
  1973 => '0',
  1974 => '0',
  1975 => '0',
  1976 => '0',
  1977 => '0',
  1978 => '0',
  1979 => '0',
  1980 => '0',
  1981 => '0',
  1982 => '0',
  1983 => '0',
  1984 => '0',
  1985 => '0',
  1986 => '0',
  1987 => '0',
  1988 => '0',
  1989 => '0',
  1990 => '0',
  1991 => '0',
  1992 => '0',
  1993 => '0',
  1994 => '0',
  1995 => '0',
  1996 => '0',
  1997 => '0',
  1998 => '0',
  1999 => '0',
  2000 => '0',
  2001 => '0',
  2002 => '0',
  2003 => '0',
  2004 => '0',
  2005 => '0',
  2006 => '0',
  2007 => '0',
  2008 => '0',
  2009 => '0',
  2010 => '0',
  2011 => '0',
  2012 => '0',
  2013 => '0',
  2014 => '0',
  2015 => '0',
  2016 => '0',
  2017 => '0',
  2018 => '0',
  2019 => '0',
  2020 => '0',
  2021 => '0',
  2022 => '0',
  2023 => '0',
  2024 => '0',
  2025 => '0',
  2026 => '0',
  2027 => '0',
  2028 => '0',
  2029 => '0',
  2030 => '0',
  2031 => '0',
  2032 => '0',
  2033 => '0',
  2034 => '0',
  2035 => '0',
  2036 => '0',
  2037 => '0',
  2038 => '0',
  2039 => '0',
  2040 => '0',
  2041 => '0',
  2042 => '0',
  2043 => '0',
  2044 => '0',
  2045 => '0',
  2046 => '0',
  2047 => '0',
  2048 => '0',
  2049 => '0',
  2050 => '0',
  2051 => '0',
  2052 => '0',
  2053 => '0',
  2054 => '0',
  2055 => '0',
  2056 => '0',
  2057 => '0',
  2058 => '0',
  2059 => '0',
  2060 => '0',
  2061 => '0',
  2062 => '0',
  2063 => '0',
  2064 => '0',
  2065 => '0',
  2066 => '0',
  2067 => '0',
  2068 => '0',
  2069 => '0',
  2070 => '0',
  2071 => '0',
  2072 => '0',
  2073 => '0',
  2074 => '0',
  2075 => '0',
  2076 => '0',
  2077 => '0',
  2078 => '0',
  2079 => '0',
  2080 => '0',
  2081 => '0',
  2082 => '0',
  2083 => '0',
  2084 => '0',
  2085 => '0',
  2086 => '0',
  2087 => '0',
  2088 => '0',
  2089 => '0',
  2090 => '0',
  2091 => '0',
  2092 => '0',
  2093 => '0',
  2094 => '0',
  2095 => '0',
  2096 => '0',
  2097 => '0',
  2098 => '0',
  2099 => '0',
  2100 => '0',
  2101 => '0',
  2102 => '0',
  2103 => '0',
  2104 => '0',
  2105 => '0',
  2106 => '0',
  2107 => '0',
  2108 => '0',
  2109 => '0',
  2110 => '0',
  2111 => '0',
  2112 => '0',
  2113 => '0',
  2114 => '0',
  2115 => '1',
  2116 => '1',
  2117 => '0',
  2118 => '0',
  2119 => '0',
  2120 => '0',
  2121 => '0',
  2122 => '0',
  2123 => '1',
  2124 => '1',
  2125 => '0',
  2126 => '0',
  2127 => '0',
  2128 => '0',
  2129 => '0',
  2130 => '0',
  2131 => '1',
  2132 => '1',
  2133 => '0',
  2134 => '0',
  2135 => '0',
  2136 => '0',
  2137 => '0',
  2138 => '0',
  2139 => '1',
  2140 => '1',
  2141 => '0',
  2142 => '0',
  2143 => '0',
  2144 => '0',
  2145 => '0',
  2146 => '0',
  2147 => '1',
  2148 => '1',
  2149 => '0',
  2150 => '0',
  2151 => '0',
  2152 => '0',
  2153 => '0',
  2154 => '0',
  2155 => '0',
  2156 => '0',
  2157 => '0',
  2158 => '0',
  2159 => '0',
  2160 => '0',
  2161 => '0',
  2162 => '0',
  2163 => '1',
  2164 => '1',
  2165 => '0',
  2166 => '0',
  2167 => '0',
  2168 => '0',
  2169 => '0',
  2170 => '0',
  2171 => '0',
  2172 => '0',
  2173 => '0',
  2174 => '0',
  2175 => '0',
  2176 => '0',
  2177 => '1',
  2178 => '1',
  2179 => '0',
  2180 => '1',
  2181 => '1',
  2182 => '0',
  2183 => '0',
  2184 => '0',
  2185 => '1',
  2186 => '1',
  2187 => '0',
  2188 => '1',
  2189 => '1',
  2190 => '0',
  2191 => '0',
  2192 => '0',
  2193 => '0',
  2194 => '0',
  2195 => '0',
  2196 => '0',
  2197 => '0',
  2198 => '0',
  2199 => '0',
  2200 => '0',
  2201 => '0',
  2202 => '0',
  2203 => '0',
  2204 => '0',
  2205 => '0',
  2206 => '0',
  2207 => '0',
  2208 => '0',
  2209 => '0',
  2210 => '0',
  2211 => '0',
  2212 => '0',
  2213 => '0',
  2214 => '0',
  2215 => '0',
  2216 => '0',
  2217 => '0',
  2218 => '0',
  2219 => '0',
  2220 => '0',
  2221 => '0',
  2222 => '0',
  2223 => '0',
  2224 => '0',
  2225 => '0',
  2226 => '0',
  2227 => '0',
  2228 => '0',
  2229 => '0',
  2230 => '0',
  2231 => '0',
  2232 => '0',
  2233 => '0',
  2234 => '0',
  2235 => '0',
  2236 => '0',
  2237 => '0',
  2238 => '0',
  2239 => '0',
  2240 => '0',
  2241 => '1',
  2242 => '1',
  2243 => '0',
  2244 => '1',
  2245 => '1',
  2246 => '0',
  2247 => '0',
  2248 => '0',
  2249 => '1',
  2250 => '1',
  2251 => '0',
  2252 => '1',
  2253 => '1',
  2254 => '0',
  2255 => '0',
  2256 => '1',
  2257 => '1',
  2258 => '1',
  2259 => '1',
  2260 => '1',
  2261 => '1',
  2262 => '1',
  2263 => '0',
  2264 => '0',
  2265 => '1',
  2266 => '1',
  2267 => '0',
  2268 => '1',
  2269 => '1',
  2270 => '0',
  2271 => '0',
  2272 => '1',
  2273 => '1',
  2274 => '1',
  2275 => '1',
  2276 => '1',
  2277 => '1',
  2278 => '1',
  2279 => '0',
  2280 => '0',
  2281 => '1',
  2282 => '1',
  2283 => '0',
  2284 => '1',
  2285 => '1',
  2286 => '0',
  2287 => '0',
  2288 => '0',
  2289 => '1',
  2290 => '1',
  2291 => '0',
  2292 => '1',
  2293 => '1',
  2294 => '0',
  2295 => '0',
  2296 => '0',
  2297 => '0',
  2298 => '0',
  2299 => '0',
  2300 => '0',
  2301 => '0',
  2302 => '0',
  2303 => '0',
  2304 => '0',
  2305 => '0',
  2306 => '0',
  2307 => '1',
  2308 => '1',
  2309 => '0',
  2310 => '0',
  2311 => '0',
  2312 => '0',
  2313 => '0',
  2314 => '1',
  2315 => '1',
  2316 => '1',
  2317 => '1',
  2318 => '1',
  2319 => '0',
  2320 => '0',
  2321 => '1',
  2322 => '1',
  2323 => '0',
  2324 => '0',
  2325 => '0',
  2326 => '0',
  2327 => '0',
  2328 => '0',
  2329 => '0',
  2330 => '1',
  2331 => '1',
  2332 => '1',
  2333 => '1',
  2334 => '0',
  2335 => '0',
  2336 => '0',
  2337 => '0',
  2338 => '0',
  2339 => '0',
  2340 => '0',
  2341 => '1',
  2342 => '1',
  2343 => '0',
  2344 => '0',
  2345 => '1',
  2346 => '1',
  2347 => '1',
  2348 => '1',
  2349 => '1',
  2350 => '0',
  2351 => '0',
  2352 => '0',
  2353 => '0',
  2354 => '0',
  2355 => '1',
  2356 => '1',
  2357 => '0',
  2358 => '0',
  2359 => '0',
  2360 => '0',
  2361 => '0',
  2362 => '0',
  2363 => '0',
  2364 => '0',
  2365 => '0',
  2366 => '0',
  2367 => '0',
  2368 => '0',
  2369 => '0',
  2370 => '0',
  2371 => '0',
  2372 => '0',
  2373 => '0',
  2374 => '0',
  2375 => '0',
  2376 => '0',
  2377 => '1',
  2378 => '1',
  2379 => '0',
  2380 => '0',
  2381 => '1',
  2382 => '1',
  2383 => '0',
  2384 => '1',
  2385 => '0',
  2386 => '1',
  2387 => '0',
  2388 => '1',
  2389 => '1',
  2390 => '0',
  2391 => '0',
  2392 => '1',
  2393 => '1',
  2394 => '0',
  2395 => '1',
  2396 => '1',
  2397 => '0',
  2398 => '0',
  2399 => '0',
  2400 => '0',
  2401 => '0',
  2402 => '1',
  2403 => '1',
  2404 => '0',
  2405 => '1',
  2406 => '1',
  2407 => '0',
  2408 => '0',
  2409 => '1',
  2410 => '1',
  2411 => '0',
  2412 => '1',
  2413 => '0',
  2414 => '1',
  2415 => '0',
  2416 => '1',
  2417 => '1',
  2418 => '0',
  2419 => '0',
  2420 => '1',
  2421 => '1',
  2422 => '0',
  2423 => '0',
  2424 => '0',
  2425 => '0',
  2426 => '0',
  2427 => '0',
  2428 => '0',
  2429 => '0',
  2430 => '0',
  2431 => '0',
  2432 => '0',
  2433 => '0',
  2434 => '1',
  2435 => '1',
  2436 => '1',
  2437 => '0',
  2438 => '0',
  2439 => '0',
  2440 => '0',
  2441 => '1',
  2442 => '1',
  2443 => '0',
  2444 => '1',
  2445 => '1',
  2446 => '0',
  2447 => '0',
  2448 => '0',
  2449 => '1',
  2450 => '1',
  2451 => '0',
  2452 => '1',
  2453 => '0',
  2454 => '0',
  2455 => '0',
  2456 => '0',
  2457 => '1',
  2458 => '1',
  2459 => '1',
  2460 => '0',
  2461 => '1',
  2462 => '1',
  2463 => '0',
  2464 => '1',
  2465 => '1',
  2466 => '0',
  2467 => '1',
  2468 => '1',
  2469 => '1',
  2470 => '0',
  2471 => '0',
  2472 => '1',
  2473 => '1',
  2474 => '0',
  2475 => '0',
  2476 => '1',
  2477 => '1',
  2478 => '1',
  2479 => '0',
  2480 => '0',
  2481 => '1',
  2482 => '1',
  2483 => '1',
  2484 => '1',
  2485 => '0',
  2486 => '1',
  2487 => '1',
  2488 => '0',
  2489 => '0',
  2490 => '0',
  2491 => '0',
  2492 => '0',
  2493 => '0',
  2494 => '0',
  2495 => '0',
  2496 => '0',
  2497 => '0',
  2498 => '0',
  2499 => '1',
  2500 => '1',
  2501 => '0',
  2502 => '0',
  2503 => '0',
  2504 => '0',
  2505 => '0',
  2506 => '0',
  2507 => '1',
  2508 => '1',
  2509 => '0',
  2510 => '0',
  2511 => '0',
  2512 => '0',
  2513 => '0',
  2514 => '1',
  2515 => '1',
  2516 => '0',
  2517 => '0',
  2518 => '0',
  2519 => '0',
  2520 => '0',
  2521 => '0',
  2522 => '0',
  2523 => '0',
  2524 => '0',
  2525 => '0',
  2526 => '0',
  2527 => '0',
  2528 => '0',
  2529 => '0',
  2530 => '0',
  2531 => '0',
  2532 => '0',
  2533 => '0',
  2534 => '0',
  2535 => '0',
  2536 => '0',
  2537 => '0',
  2538 => '0',
  2539 => '0',
  2540 => '0',
  2541 => '0',
  2542 => '0',
  2543 => '0',
  2544 => '0',
  2545 => '0',
  2546 => '0',
  2547 => '0',
  2548 => '0',
  2549 => '0',
  2550 => '0',
  2551 => '0',
  2552 => '0',
  2553 => '0',
  2554 => '0',
  2555 => '0',
  2556 => '0',
  2557 => '0',
  2558 => '0',
  2559 => '0',
  2560 => '0',
  2561 => '0',
  2562 => '0',
  2563 => '0',
  2564 => '1',
  2565 => '1',
  2566 => '0',
  2567 => '0',
  2568 => '0',
  2569 => '0',
  2570 => '0',
  2571 => '1',
  2572 => '1',
  2573 => '0',
  2574 => '0',
  2575 => '0',
  2576 => '0',
  2577 => '0',
  2578 => '1',
  2579 => '1',
  2580 => '0',
  2581 => '0',
  2582 => '0',
  2583 => '0',
  2584 => '0',
  2585 => '0',
  2586 => '1',
  2587 => '1',
  2588 => '0',
  2589 => '0',
  2590 => '0',
  2591 => '0',
  2592 => '0',
  2593 => '0',
  2594 => '1',
  2595 => '1',
  2596 => '0',
  2597 => '0',
  2598 => '0',
  2599 => '0',
  2600 => '0',
  2601 => '0',
  2602 => '0',
  2603 => '1',
  2604 => '1',
  2605 => '0',
  2606 => '0',
  2607 => '0',
  2608 => '0',
  2609 => '0',
  2610 => '0',
  2611 => '0',
  2612 => '1',
  2613 => '1',
  2614 => '0',
  2615 => '0',
  2616 => '0',
  2617 => '0',
  2618 => '0',
  2619 => '0',
  2620 => '0',
  2621 => '0',
  2622 => '0',
  2623 => '0',
  2624 => '0',
  2625 => '0',
  2626 => '1',
  2627 => '1',
  2628 => '0',
  2629 => '0',
  2630 => '0',
  2631 => '0',
  2632 => '0',
  2633 => '0',
  2634 => '0',
  2635 => '1',
  2636 => '1',
  2637 => '0',
  2638 => '0',
  2639 => '0',
  2640 => '0',
  2641 => '0',
  2642 => '0',
  2643 => '0',
  2644 => '1',
  2645 => '1',
  2646 => '0',
  2647 => '0',
  2648 => '0',
  2649 => '0',
  2650 => '0',
  2651 => '0',
  2652 => '1',
  2653 => '1',
  2654 => '0',
  2655 => '0',
  2656 => '0',
  2657 => '0',
  2658 => '0',
  2659 => '0',
  2660 => '1',
  2661 => '1',
  2662 => '0',
  2663 => '0',
  2664 => '0',
  2665 => '0',
  2666 => '0',
  2667 => '1',
  2668 => '1',
  2669 => '0',
  2670 => '0',
  2671 => '0',
  2672 => '0',
  2673 => '0',
  2674 => '1',
  2675 => '1',
  2676 => '0',
  2677 => '0',
  2678 => '0',
  2679 => '0',
  2680 => '0',
  2681 => '0',
  2682 => '0',
  2683 => '0',
  2684 => '0',
  2685 => '0',
  2686 => '0',
  2687 => '0',
  2688 => '0',
  2689 => '0',
  2690 => '0',
  2691 => '0',
  2692 => '0',
  2693 => '0',
  2694 => '0',
  2695 => '0',
  2696 => '0',
  2697 => '1',
  2698 => '1',
  2699 => '0',
  2700 => '0',
  2701 => '1',
  2702 => '1',
  2703 => '0',
  2704 => '0',
  2705 => '0',
  2706 => '1',
  2707 => '1',
  2708 => '1',
  2709 => '1',
  2710 => '0',
  2711 => '0',
  2712 => '1',
  2713 => '1',
  2714 => '1',
  2715 => '1',
  2716 => '1',
  2717 => '1',
  2718 => '1',
  2719 => '1',
  2720 => '0',
  2721 => '0',
  2722 => '1',
  2723 => '1',
  2724 => '1',
  2725 => '1',
  2726 => '0',
  2727 => '0',
  2728 => '0',
  2729 => '1',
  2730 => '1',
  2731 => '0',
  2732 => '0',
  2733 => '1',
  2734 => '1',
  2735 => '0',
  2736 => '0',
  2737 => '0',
  2738 => '0',
  2739 => '0',
  2740 => '0',
  2741 => '0',
  2742 => '0',
  2743 => '0',
  2744 => '0',
  2745 => '0',
  2746 => '0',
  2747 => '0',
  2748 => '0',
  2749 => '0',
  2750 => '0',
  2751 => '0',
  2752 => '0',
  2753 => '0',
  2754 => '0',
  2755 => '0',
  2756 => '0',
  2757 => '0',
  2758 => '0',
  2759 => '0',
  2760 => '0',
  2761 => '0',
  2762 => '0',
  2763 => '1',
  2764 => '1',
  2765 => '0',
  2766 => '0',
  2767 => '0',
  2768 => '0',
  2769 => '0',
  2770 => '0',
  2771 => '1',
  2772 => '1',
  2773 => '0',
  2774 => '0',
  2775 => '0',
  2776 => '0',
  2777 => '1',
  2778 => '1',
  2779 => '1',
  2780 => '1',
  2781 => '1',
  2782 => '1',
  2783 => '0',
  2784 => '0',
  2785 => '0',
  2786 => '0',
  2787 => '1',
  2788 => '1',
  2789 => '0',
  2790 => '0',
  2791 => '0',
  2792 => '0',
  2793 => '0',
  2794 => '0',
  2795 => '1',
  2796 => '1',
  2797 => '0',
  2798 => '0',
  2799 => '0',
  2800 => '0',
  2801 => '0',
  2802 => '0',
  2803 => '0',
  2804 => '0',
  2805 => '0',
  2806 => '0',
  2807 => '0',
  2808 => '0',
  2809 => '0',
  2810 => '0',
  2811 => '0',
  2812 => '0',
  2813 => '0',
  2814 => '0',
  2815 => '0',
  2816 => '0',
  2817 => '0',
  2818 => '0',
  2819 => '0',
  2820 => '0',
  2821 => '0',
  2822 => '0',
  2823 => '0',
  2824 => '0',
  2825 => '0',
  2826 => '0',
  2827 => '0',
  2828 => '0',
  2829 => '0',
  2830 => '0',
  2831 => '0',
  2832 => '0',
  2833 => '0',
  2834 => '0',
  2835 => '0',
  2836 => '0',
  2837 => '0',
  2838 => '0',
  2839 => '0',
  2840 => '0',
  2841 => '0',
  2842 => '0',
  2843 => '0',
  2844 => '0',
  2845 => '0',
  2846 => '0',
  2847 => '0',
  2848 => '0',
  2849 => '0',
  2850 => '0',
  2851 => '0',
  2852 => '0',
  2853 => '0',
  2854 => '0',
  2855 => '0',
  2856 => '0',
  2857 => '0',
  2858 => '0',
  2859 => '1',
  2860 => '1',
  2861 => '0',
  2862 => '0',
  2863 => '0',
  2864 => '0',
  2865 => '0',
  2866 => '0',
  2867 => '1',
  2868 => '1',
  2869 => '0',
  2870 => '0',
  2871 => '0',
  2872 => '0',
  2873 => '0',
  2874 => '1',
  2875 => '1',
  2876 => '0',
  2877 => '0',
  2878 => '0',
  2879 => '0',
  2880 => '0',
  2881 => '0',
  2882 => '0',
  2883 => '0',
  2884 => '0',
  2885 => '0',
  2886 => '0',
  2887 => '0',
  2888 => '0',
  2889 => '0',
  2890 => '0',
  2891 => '0',
  2892 => '0',
  2893 => '0',
  2894 => '0',
  2895 => '0',
  2896 => '0',
  2897 => '0',
  2898 => '0',
  2899 => '0',
  2900 => '0',
  2901 => '0',
  2902 => '0',
  2903 => '0',
  2904 => '0',
  2905 => '1',
  2906 => '1',
  2907 => '1',
  2908 => '1',
  2909 => '1',
  2910 => '1',
  2911 => '0',
  2912 => '0',
  2913 => '0',
  2914 => '0',
  2915 => '0',
  2916 => '0',
  2917 => '0',
  2918 => '0',
  2919 => '0',
  2920 => '0',
  2921 => '0',
  2922 => '0',
  2923 => '0',
  2924 => '0',
  2925 => '0',
  2926 => '0',
  2927 => '0',
  2928 => '0',
  2929 => '0',
  2930 => '0',
  2931 => '0',
  2932 => '0',
  2933 => '0',
  2934 => '0',
  2935 => '0',
  2936 => '0',
  2937 => '0',
  2938 => '0',
  2939 => '0',
  2940 => '0',
  2941 => '0',
  2942 => '0',
  2943 => '0',
  2944 => '0',
  2945 => '0',
  2946 => '0',
  2947 => '0',
  2948 => '0',
  2949 => '0',
  2950 => '0',
  2951 => '0',
  2952 => '0',
  2953 => '0',
  2954 => '0',
  2955 => '0',
  2956 => '0',
  2957 => '0',
  2958 => '0',
  2959 => '0',
  2960 => '0',
  2961 => '0',
  2962 => '0',
  2963 => '0',
  2964 => '0',
  2965 => '0',
  2966 => '0',
  2967 => '0',
  2968 => '0',
  2969 => '0',
  2970 => '0',
  2971 => '0',
  2972 => '0',
  2973 => '0',
  2974 => '0',
  2975 => '0',
  2976 => '0',
  2977 => '0',
  2978 => '0',
  2979 => '0',
  2980 => '0',
  2981 => '0',
  2982 => '0',
  2983 => '0',
  2984 => '0',
  2985 => '0',
  2986 => '0',
  2987 => '1',
  2988 => '1',
  2989 => '0',
  2990 => '0',
  2991 => '0',
  2992 => '0',
  2993 => '0',
  2994 => '0',
  2995 => '1',
  2996 => '1',
  2997 => '0',
  2998 => '0',
  2999 => '0',
  3000 => '0',
  3001 => '0',
  3002 => '0',
  3003 => '0',
  3004 => '0',
  3005 => '0',
  3006 => '0',
  3007 => '0',
  3008 => '0',
  3009 => '0',
  3010 => '0',
  3011 => '0',
  3012 => '0',
  3013 => '0',
  3014 => '1',
  3015 => '1',
  3016 => '0',
  3017 => '0',
  3018 => '0',
  3019 => '0',
  3020 => '0',
  3021 => '1',
  3022 => '1',
  3023 => '0',
  3024 => '0',
  3025 => '0',
  3026 => '0',
  3027 => '0',
  3028 => '1',
  3029 => '1',
  3030 => '0',
  3031 => '0',
  3032 => '0',
  3033 => '0',
  3034 => '0',
  3035 => '1',
  3036 => '1',
  3037 => '0',
  3038 => '0',
  3039 => '0',
  3040 => '0',
  3041 => '0',
  3042 => '1',
  3043 => '1',
  3044 => '0',
  3045 => '0',
  3046 => '0',
  3047 => '0',
  3048 => '0',
  3049 => '1',
  3050 => '1',
  3051 => '0',
  3052 => '0',
  3053 => '0',
  3054 => '0',
  3055 => '0',
  3056 => '1',
  3057 => '1',
  3058 => '0',
  3059 => '0',
  3060 => '0',
  3061 => '0',
  3062 => '0',
  3063 => '0',
  3064 => '0',
  3065 => '0',
  3066 => '0',
  3067 => '0',
  3068 => '0',
  3069 => '0',
  3070 => '0',
  3071 => '0',
  3072 => '0',
  3073 => '0',
  3074 => '1',
  3075 => '1',
  3076 => '1',
  3077 => '1',
  3078 => '0',
  3079 => '0',
  3080 => '0',
  3081 => '1',
  3082 => '1',
  3083 => '0',
  3084 => '0',
  3085 => '1',
  3086 => '1',
  3087 => '0',
  3088 => '0',
  3089 => '1',
  3090 => '1',
  3091 => '0',
  3092 => '1',
  3093 => '1',
  3094 => '1',
  3095 => '0',
  3096 => '0',
  3097 => '1',
  3098 => '1',
  3099 => '1',
  3100 => '1',
  3101 => '1',
  3102 => '1',
  3103 => '0',
  3104 => '0',
  3105 => '1',
  3106 => '1',
  3107 => '1',
  3108 => '0',
  3109 => '1',
  3110 => '1',
  3111 => '0',
  3112 => '0',
  3113 => '1',
  3114 => '1',
  3115 => '0',
  3116 => '0',
  3117 => '1',
  3118 => '1',
  3119 => '0',
  3120 => '0',
  3121 => '0',
  3122 => '1',
  3123 => '1',
  3124 => '1',
  3125 => '1',
  3126 => '0',
  3127 => '0',
  3128 => '0',
  3129 => '0',
  3130 => '0',
  3131 => '0',
  3132 => '0',
  3133 => '0',
  3134 => '0',
  3135 => '0',
  3136 => '0',
  3137 => '0',
  3138 => '0',
  3139 => '1',
  3140 => '1',
  3141 => '0',
  3142 => '0',
  3143 => '0',
  3144 => '0',
  3145 => '0',
  3146 => '1',
  3147 => '1',
  3148 => '1',
  3149 => '0',
  3150 => '0',
  3151 => '0',
  3152 => '0',
  3153 => '1',
  3154 => '1',
  3155 => '1',
  3156 => '1',
  3157 => '0',
  3158 => '0',
  3159 => '0',
  3160 => '0',
  3161 => '0',
  3162 => '0',
  3163 => '1',
  3164 => '1',
  3165 => '0',
  3166 => '0',
  3167 => '0',
  3168 => '0',
  3169 => '0',
  3170 => '0',
  3171 => '1',
  3172 => '1',
  3173 => '0',
  3174 => '0',
  3175 => '0',
  3176 => '0',
  3177 => '0',
  3178 => '0',
  3179 => '1',
  3180 => '1',
  3181 => '0',
  3182 => '0',
  3183 => '0',
  3184 => '0',
  3185 => '0',
  3186 => '0',
  3187 => '1',
  3188 => '1',
  3189 => '0',
  3190 => '0',
  3191 => '0',
  3192 => '0',
  3193 => '0',
  3194 => '0',
  3195 => '0',
  3196 => '0',
  3197 => '0',
  3198 => '0',
  3199 => '0',
  3200 => '0',
  3201 => '0',
  3202 => '1',
  3203 => '1',
  3204 => '1',
  3205 => '1',
  3206 => '0',
  3207 => '0',
  3208 => '0',
  3209 => '1',
  3210 => '1',
  3211 => '0',
  3212 => '0',
  3213 => '1',
  3214 => '1',
  3215 => '0',
  3216 => '0',
  3217 => '0',
  3218 => '0',
  3219 => '0',
  3220 => '0',
  3221 => '1',
  3222 => '1',
  3223 => '0',
  3224 => '0',
  3225 => '0',
  3226 => '0',
  3227 => '0',
  3228 => '1',
  3229 => '1',
  3230 => '0',
  3231 => '0',
  3232 => '0',
  3233 => '0',
  3234 => '0',
  3235 => '1',
  3236 => '1',
  3237 => '0',
  3238 => '0',
  3239 => '0',
  3240 => '0',
  3241 => '0',
  3242 => '1',
  3243 => '1',
  3244 => '0',
  3245 => '0',
  3246 => '0',
  3247 => '0',
  3248 => '0',
  3249 => '1',
  3250 => '1',
  3251 => '1',
  3252 => '1',
  3253 => '1',
  3254 => '1',
  3255 => '0',
  3256 => '0',
  3257 => '0',
  3258 => '0',
  3259 => '0',
  3260 => '0',
  3261 => '0',
  3262 => '0',
  3263 => '0',
  3264 => '0',
  3265 => '0',
  3266 => '1',
  3267 => '1',
  3268 => '1',
  3269 => '1',
  3270 => '0',
  3271 => '0',
  3272 => '0',
  3273 => '1',
  3274 => '1',
  3275 => '0',
  3276 => '0',
  3277 => '1',
  3278 => '1',
  3279 => '0',
  3280 => '0',
  3281 => '0',
  3282 => '0',
  3283 => '0',
  3284 => '0',
  3285 => '1',
  3286 => '1',
  3287 => '0',
  3288 => '0',
  3289 => '0',
  3290 => '0',
  3291 => '1',
  3292 => '1',
  3293 => '1',
  3294 => '0',
  3295 => '0',
  3296 => '0',
  3297 => '0',
  3298 => '0',
  3299 => '0',
  3300 => '0',
  3301 => '1',
  3302 => '1',
  3303 => '0',
  3304 => '0',
  3305 => '1',
  3306 => '1',
  3307 => '0',
  3308 => '0',
  3309 => '1',
  3310 => '1',
  3311 => '0',
  3312 => '0',
  3313 => '0',
  3314 => '1',
  3315 => '1',
  3316 => '1',
  3317 => '1',
  3318 => '0',
  3319 => '0',
  3320 => '0',
  3321 => '0',
  3322 => '0',
  3323 => '0',
  3324 => '0',
  3325 => '0',
  3326 => '0',
  3327 => '0',
  3328 => '0',
  3329 => '0',
  3330 => '0',
  3331 => '1',
  3332 => '1',
  3333 => '1',
  3334 => '0',
  3335 => '0',
  3336 => '0',
  3337 => '0',
  3338 => '1',
  3339 => '1',
  3340 => '1',
  3341 => '1',
  3342 => '0',
  3343 => '0',
  3344 => '0',
  3345 => '1',
  3346 => '1',
  3347 => '0',
  3348 => '1',
  3349 => '1',
  3350 => '0',
  3351 => '0',
  3352 => '1',
  3353 => '1',
  3354 => '0',
  3355 => '0',
  3356 => '1',
  3357 => '1',
  3358 => '0',
  3359 => '0',
  3360 => '1',
  3361 => '1',
  3362 => '1',
  3363 => '1',
  3364 => '1',
  3365 => '1',
  3366 => '1',
  3367 => '0',
  3368 => '0',
  3369 => '0',
  3370 => '0',
  3371 => '0',
  3372 => '1',
  3373 => '1',
  3374 => '0',
  3375 => '0',
  3376 => '0',
  3377 => '0',
  3378 => '0',
  3379 => '0',
  3380 => '1',
  3381 => '1',
  3382 => '0',
  3383 => '0',
  3384 => '0',
  3385 => '0',
  3386 => '0',
  3387 => '0',
  3388 => '0',
  3389 => '0',
  3390 => '0',
  3391 => '0',
  3392 => '0',
  3393 => '1',
  3394 => '1',
  3395 => '1',
  3396 => '1',
  3397 => '1',
  3398 => '1',
  3399 => '0',
  3400 => '0',
  3401 => '1',
  3402 => '1',
  3403 => '0',
  3404 => '0',
  3405 => '0',
  3406 => '0',
  3407 => '0',
  3408 => '0',
  3409 => '1',
  3410 => '1',
  3411 => '1',
  3412 => '1',
  3413 => '1',
  3414 => '0',
  3415 => '0',
  3416 => '0',
  3417 => '0',
  3418 => '0',
  3419 => '0',
  3420 => '0',
  3421 => '1',
  3422 => '1',
  3423 => '0',
  3424 => '0',
  3425 => '0',
  3426 => '0',
  3427 => '0',
  3428 => '0',
  3429 => '1',
  3430 => '1',
  3431 => '0',
  3432 => '0',
  3433 => '1',
  3434 => '1',
  3435 => '0',
  3436 => '0',
  3437 => '1',
  3438 => '1',
  3439 => '0',
  3440 => '0',
  3441 => '0',
  3442 => '1',
  3443 => '1',
  3444 => '1',
  3445 => '1',
  3446 => '0',
  3447 => '0',
  3448 => '0',
  3449 => '0',
  3450 => '0',
  3451 => '0',
  3452 => '0',
  3453 => '0',
  3454 => '0',
  3455 => '0',
  3456 => '0',
  3457 => '0',
  3458 => '0',
  3459 => '1',
  3460 => '1',
  3461 => '1',
  3462 => '0',
  3463 => '0',
  3464 => '0',
  3465 => '0',
  3466 => '1',
  3467 => '1',
  3468 => '0',
  3469 => '0',
  3470 => '0',
  3471 => '0',
  3472 => '0',
  3473 => '1',
  3474 => '1',
  3475 => '0',
  3476 => '0',
  3477 => '0',
  3478 => '0',
  3479 => '0',
  3480 => '0',
  3481 => '1',
  3482 => '1',
  3483 => '1',
  3484 => '1',
  3485 => '1',
  3486 => '0',
  3487 => '0',
  3488 => '0',
  3489 => '1',
  3490 => '1',
  3491 => '0',
  3492 => '0',
  3493 => '1',
  3494 => '1',
  3495 => '0',
  3496 => '0',
  3497 => '1',
  3498 => '1',
  3499 => '0',
  3500 => '0',
  3501 => '1',
  3502 => '1',
  3503 => '0',
  3504 => '0',
  3505 => '0',
  3506 => '1',
  3507 => '1',
  3508 => '1',
  3509 => '1',
  3510 => '0',
  3511 => '0',
  3512 => '0',
  3513 => '0',
  3514 => '0',
  3515 => '0',
  3516 => '0',
  3517 => '0',
  3518 => '0',
  3519 => '0',
  3520 => '0',
  3521 => '1',
  3522 => '1',
  3523 => '1',
  3524 => '1',
  3525 => '1',
  3526 => '1',
  3527 => '0',
  3528 => '0',
  3529 => '0',
  3530 => '0',
  3531 => '0',
  3532 => '0',
  3533 => '1',
  3534 => '1',
  3535 => '0',
  3536 => '0',
  3537 => '0',
  3538 => '0',
  3539 => '0',
  3540 => '0',
  3541 => '1',
  3542 => '1',
  3543 => '0',
  3544 => '0',
  3545 => '0',
  3546 => '0',
  3547 => '0',
  3548 => '1',
  3549 => '1',
  3550 => '0',
  3551 => '0',
  3552 => '0',
  3553 => '0',
  3554 => '0',
  3555 => '1',
  3556 => '1',
  3557 => '0',
  3558 => '0',
  3559 => '0',
  3560 => '0',
  3561 => '0',
  3562 => '0',
  3563 => '1',
  3564 => '1',
  3565 => '0',
  3566 => '0',
  3567 => '0',
  3568 => '0',
  3569 => '0',
  3570 => '0',
  3571 => '1',
  3572 => '1',
  3573 => '0',
  3574 => '0',
  3575 => '0',
  3576 => '0',
  3577 => '0',
  3578 => '0',
  3579 => '0',
  3580 => '0',
  3581 => '0',
  3582 => '0',
  3583 => '0',
  3584 => '0',
  3585 => '0',
  3586 => '1',
  3587 => '1',
  3588 => '1',
  3589 => '1',
  3590 => '0',
  3591 => '0',
  3592 => '0',
  3593 => '1',
  3594 => '1',
  3595 => '0',
  3596 => '0',
  3597 => '1',
  3598 => '1',
  3599 => '0',
  3600 => '0',
  3601 => '1',
  3602 => '1',
  3603 => '0',
  3604 => '0',
  3605 => '1',
  3606 => '1',
  3607 => '0',
  3608 => '0',
  3609 => '0',
  3610 => '1',
  3611 => '1',
  3612 => '1',
  3613 => '1',
  3614 => '0',
  3615 => '0',
  3616 => '0',
  3617 => '1',
  3618 => '1',
  3619 => '0',
  3620 => '0',
  3621 => '1',
  3622 => '1',
  3623 => '0',
  3624 => '0',
  3625 => '1',
  3626 => '1',
  3627 => '0',
  3628 => '0',
  3629 => '1',
  3630 => '1',
  3631 => '0',
  3632 => '0',
  3633 => '0',
  3634 => '1',
  3635 => '1',
  3636 => '1',
  3637 => '1',
  3638 => '0',
  3639 => '0',
  3640 => '0',
  3641 => '0',
  3642 => '0',
  3643 => '0',
  3644 => '0',
  3645 => '0',
  3646 => '0',
  3647 => '0',
  3648 => '0',
  3649 => '0',
  3650 => '1',
  3651 => '1',
  3652 => '1',
  3653 => '1',
  3654 => '0',
  3655 => '0',
  3656 => '0',
  3657 => '1',
  3658 => '1',
  3659 => '0',
  3660 => '0',
  3661 => '1',
  3662 => '1',
  3663 => '0',
  3664 => '0',
  3665 => '1',
  3666 => '1',
  3667 => '0',
  3668 => '0',
  3669 => '1',
  3670 => '1',
  3671 => '0',
  3672 => '0',
  3673 => '0',
  3674 => '1',
  3675 => '1',
  3676 => '1',
  3677 => '1',
  3678 => '1',
  3679 => '0',
  3680 => '0',
  3681 => '0',
  3682 => '0',
  3683 => '0',
  3684 => '0',
  3685 => '1',
  3686 => '1',
  3687 => '0',
  3688 => '0',
  3689 => '0',
  3690 => '0',
  3691 => '0',
  3692 => '1',
  3693 => '1',
  3694 => '0',
  3695 => '0',
  3696 => '0',
  3697 => '0',
  3698 => '1',
  3699 => '1',
  3700 => '1',
  3701 => '0',
  3702 => '0',
  3703 => '0',
  3704 => '0',
  3705 => '0',
  3706 => '0',
  3707 => '0',
  3708 => '0',
  3709 => '0',
  3710 => '0',
  3711 => '0',
  3712 => '0',
  3713 => '0',
  3714 => '0',
  3715 => '0',
  3716 => '0',
  3717 => '0',
  3718 => '0',
  3719 => '0',
  3720 => '0',
  3721 => '0',
  3722 => '0',
  3723 => '1',
  3724 => '1',
  3725 => '0',
  3726 => '0',
  3727 => '0',
  3728 => '0',
  3729 => '0',
  3730 => '0',
  3731 => '1',
  3732 => '1',
  3733 => '0',
  3734 => '0',
  3735 => '0',
  3736 => '0',
  3737 => '0',
  3738 => '0',
  3739 => '0',
  3740 => '0',
  3741 => '0',
  3742 => '0',
  3743 => '0',
  3744 => '0',
  3745 => '0',
  3746 => '0',
  3747 => '0',
  3748 => '0',
  3749 => '0',
  3750 => '0',
  3751 => '0',
  3752 => '0',
  3753 => '0',
  3754 => '0',
  3755 => '1',
  3756 => '1',
  3757 => '0',
  3758 => '0',
  3759 => '0',
  3760 => '0',
  3761 => '0',
  3762 => '0',
  3763 => '1',
  3764 => '1',
  3765 => '0',
  3766 => '0',
  3767 => '0',
  3768 => '0',
  3769 => '0',
  3770 => '0',
  3771 => '0',
  3772 => '0',
  3773 => '0',
  3774 => '0',
  3775 => '0',
  3776 => '0',
  3777 => '0',
  3778 => '0',
  3779 => '0',
  3780 => '0',
  3781 => '0',
  3782 => '0',
  3783 => '0',
  3784 => '0',
  3785 => '0',
  3786 => '0',
  3787 => '1',
  3788 => '1',
  3789 => '0',
  3790 => '0',
  3791 => '0',
  3792 => '0',
  3793 => '0',
  3794 => '0',
  3795 => '1',
  3796 => '1',
  3797 => '0',
  3798 => '0',
  3799 => '0',
  3800 => '0',
  3801 => '0',
  3802 => '0',
  3803 => '0',
  3804 => '0',
  3805 => '0',
  3806 => '0',
  3807 => '0',
  3808 => '0',
  3809 => '0',
  3810 => '0',
  3811 => '0',
  3812 => '0',
  3813 => '0',
  3814 => '0',
  3815 => '0',
  3816 => '0',
  3817 => '0',
  3818 => '0',
  3819 => '1',
  3820 => '1',
  3821 => '0',
  3822 => '0',
  3823 => '0',
  3824 => '0',
  3825 => '0',
  3826 => '0',
  3827 => '1',
  3828 => '1',
  3829 => '0',
  3830 => '0',
  3831 => '0',
  3832 => '0',
  3833 => '0',
  3834 => '1',
  3835 => '1',
  3836 => '0',
  3837 => '0',
  3838 => '0',
  3839 => '0',
  3840 => '0',
  3841 => '0',
  3842 => '0',
  3843 => '0',
  3844 => '0',
  3845 => '0',
  3846 => '0',
  3847 => '0',
  3848 => '0',
  3849 => '0',
  3850 => '0',
  3851 => '0',
  3852 => '0',
  3853 => '1',
  3854 => '1',
  3855 => '0',
  3856 => '0',
  3857 => '0',
  3858 => '0',
  3859 => '1',
  3860 => '1',
  3861 => '0',
  3862 => '0',
  3863 => '0',
  3864 => '0',
  3865 => '1',
  3866 => '1',
  3867 => '0',
  3868 => '0',
  3869 => '0',
  3870 => '0',
  3871 => '0',
  3872 => '0',
  3873 => '0',
  3874 => '0',
  3875 => '1',
  3876 => '1',
  3877 => '0',
  3878 => '0',
  3879 => '0',
  3880 => '0',
  3881 => '0',
  3882 => '0',
  3883 => '0',
  3884 => '0',
  3885 => '1',
  3886 => '1',
  3887 => '0',
  3888 => '0',
  3889 => '0',
  3890 => '0',
  3891 => '0',
  3892 => '0',
  3893 => '0',
  3894 => '0',
  3895 => '0',
  3896 => '0',
  3897 => '0',
  3898 => '0',
  3899 => '0',
  3900 => '0',
  3901 => '0',
  3902 => '0',
  3903 => '0',
  3904 => '0',
  3905 => '0',
  3906 => '0',
  3907 => '0',
  3908 => '0',
  3909 => '0',
  3910 => '0',
  3911 => '0',
  3912 => '0',
  3913 => '0',
  3914 => '0',
  3915 => '0',
  3916 => '0',
  3917 => '0',
  3918 => '0',
  3919 => '0',
  3920 => '0',
  3921 => '1',
  3922 => '1',
  3923 => '1',
  3924 => '1',
  3925 => '1',
  3926 => '1',
  3927 => '0',
  3928 => '0',
  3929 => '0',
  3930 => '0',
  3931 => '0',
  3932 => '0',
  3933 => '0',
  3934 => '0',
  3935 => '0',
  3936 => '0',
  3937 => '1',
  3938 => '1',
  3939 => '1',
  3940 => '1',
  3941 => '1',
  3942 => '1',
  3943 => '0',
  3944 => '0',
  3945 => '0',
  3946 => '0',
  3947 => '0',
  3948 => '0',
  3949 => '0',
  3950 => '0',
  3951 => '0',
  3952 => '0',
  3953 => '0',
  3954 => '0',
  3955 => '0',
  3956 => '0',
  3957 => '0',
  3958 => '0',
  3959 => '0',
  3960 => '0',
  3961 => '0',
  3962 => '0',
  3963 => '0',
  3964 => '0',
  3965 => '0',
  3966 => '0',
  3967 => '0',
  3968 => '0',
  3969 => '0',
  3970 => '0',
  3971 => '0',
  3972 => '0',
  3973 => '0',
  3974 => '0',
  3975 => '0',
  3976 => '0',
  3977 => '1',
  3978 => '1',
  3979 => '0',
  3980 => '0',
  3981 => '0',
  3982 => '0',
  3983 => '0',
  3984 => '0',
  3985 => '0',
  3986 => '0',
  3987 => '1',
  3988 => '1',
  3989 => '0',
  3990 => '0',
  3991 => '0',
  3992 => '0',
  3993 => '0',
  3994 => '0',
  3995 => '0',
  3996 => '0',
  3997 => '1',
  3998 => '1',
  3999 => '0',
  4000 => '0',
  4001 => '0',
  4002 => '0',
  4003 => '1',
  4004 => '1',
  4005 => '0',
  4006 => '0',
  4007 => '0',
  4008 => '0',
  4009 => '1',
  4010 => '1',
  4011 => '0',
  4012 => '0',
  4013 => '0',
  4014 => '0',
  4015 => '0',
  4016 => '0',
  4017 => '0',
  4018 => '0',
  4019 => '0',
  4020 => '0',
  4021 => '0',
  4022 => '0',
  4023 => '0',
  4024 => '0',
  4025 => '0',
  4026 => '0',
  4027 => '0',
  4028 => '0',
  4029 => '0',
  4030 => '0',
  4031 => '0',
  4032 => '0',
  4033 => '0',
  4034 => '1',
  4035 => '1',
  4036 => '1',
  4037 => '1',
  4038 => '0',
  4039 => '0',
  4040 => '0',
  4041 => '1',
  4042 => '1',
  4043 => '0',
  4044 => '0',
  4045 => '1',
  4046 => '1',
  4047 => '0',
  4048 => '0',
  4049 => '0',
  4050 => '0',
  4051 => '0',
  4052 => '0',
  4053 => '1',
  4054 => '1',
  4055 => '0',
  4056 => '0',
  4057 => '0',
  4058 => '0',
  4059 => '0',
  4060 => '1',
  4061 => '1',
  4062 => '0',
  4063 => '0',
  4064 => '0',
  4065 => '0',
  4066 => '0',
  4067 => '1',
  4068 => '1',
  4069 => '0',
  4070 => '0',
  4071 => '0',
  4072 => '0',
  4073 => '0',
  4074 => '0',
  4075 => '0',
  4076 => '0',
  4077 => '0',
  4078 => '0',
  4079 => '0',
  4080 => '0',
  4081 => '0',
  4082 => '0',
  4083 => '1',
  4084 => '1',
  4085 => '0',
  4086 => '0',
  4087 => '0',
  4088 => '0',
  4089 => '0',
  4090 => '0',
  4091 => '0',
  4092 => '0',
  4093 => '0',
  4094 => '0',
  4095 => '0',
  4096 => '0',
  4097 => '1',
  4098 => '1',
  4099 => '1',
  4100 => '1',
  4101 => '1',
  4102 => '0',
  4103 => '0',
  4104 => '1',
  4105 => '1',
  4106 => '0',
  4107 => '0',
  4108 => '0',
  4109 => '1',
  4110 => '1',
  4111 => '0',
  4112 => '1',
  4113 => '1',
  4114 => '0',
  4115 => '1',
  4116 => '1',
  4117 => '1',
  4118 => '1',
  4119 => '0',
  4120 => '1',
  4121 => '1',
  4122 => '0',
  4123 => '1',
  4124 => '0',
  4125 => '1',
  4126 => '1',
  4127 => '0',
  4128 => '1',
  4129 => '1',
  4130 => '0',
  4131 => '1',
  4132 => '1',
  4133 => '1',
  4134 => '1',
  4135 => '0',
  4136 => '1',
  4137 => '1',
  4138 => '0',
  4139 => '0',
  4140 => '0',
  4141 => '0',
  4142 => '0',
  4143 => '0',
  4144 => '0',
  4145 => '1',
  4146 => '1',
  4147 => '1',
  4148 => '1',
  4149 => '0',
  4150 => '0',
  4151 => '0',
  4152 => '0',
  4153 => '0',
  4154 => '0',
  4155 => '0',
  4156 => '0',
  4157 => '0',
  4158 => '0',
  4159 => '0',
  4160 => '0',
  4161 => '0',
  4162 => '1',
  4163 => '1',
  4164 => '1',
  4165 => '1',
  4166 => '0',
  4167 => '0',
  4168 => '0',
  4169 => '1',
  4170 => '1',
  4171 => '0',
  4172 => '0',
  4173 => '1',
  4174 => '1',
  4175 => '0',
  4176 => '0',
  4177 => '1',
  4178 => '1',
  4179 => '0',
  4180 => '0',
  4181 => '1',
  4182 => '1',
  4183 => '0',
  4184 => '0',
  4185 => '1',
  4186 => '1',
  4187 => '1',
  4188 => '1',
  4189 => '1',
  4190 => '1',
  4191 => '0',
  4192 => '0',
  4193 => '1',
  4194 => '1',
  4195 => '0',
  4196 => '0',
  4197 => '1',
  4198 => '1',
  4199 => '0',
  4200 => '0',
  4201 => '1',
  4202 => '1',
  4203 => '0',
  4204 => '0',
  4205 => '1',
  4206 => '1',
  4207 => '0',
  4208 => '0',
  4209 => '1',
  4210 => '1',
  4211 => '0',
  4212 => '0',
  4213 => '1',
  4214 => '1',
  4215 => '0',
  4216 => '0',
  4217 => '0',
  4218 => '0',
  4219 => '0',
  4220 => '0',
  4221 => '0',
  4222 => '0',
  4223 => '0',
  4224 => '0',
  4225 => '1',
  4226 => '1',
  4227 => '1',
  4228 => '1',
  4229 => '1',
  4230 => '0',
  4231 => '0',
  4232 => '0',
  4233 => '1',
  4234 => '1',
  4235 => '0',
  4236 => '0',
  4237 => '1',
  4238 => '1',
  4239 => '0',
  4240 => '0',
  4241 => '1',
  4242 => '1',
  4243 => '0',
  4244 => '0',
  4245 => '1',
  4246 => '1',
  4247 => '0',
  4248 => '0',
  4249 => '1',
  4250 => '1',
  4251 => '1',
  4252 => '1',
  4253 => '1',
  4254 => '0',
  4255 => '0',
  4256 => '0',
  4257 => '1',
  4258 => '1',
  4259 => '0',
  4260 => '0',
  4261 => '1',
  4262 => '1',
  4263 => '0',
  4264 => '0',
  4265 => '1',
  4266 => '1',
  4267 => '0',
  4268 => '0',
  4269 => '1',
  4270 => '1',
  4271 => '0',
  4272 => '0',
  4273 => '1',
  4274 => '1',
  4275 => '1',
  4276 => '1',
  4277 => '1',
  4278 => '0',
  4279 => '0',
  4280 => '0',
  4281 => '0',
  4282 => '0',
  4283 => '0',
  4284 => '0',
  4285 => '0',
  4286 => '0',
  4287 => '0',
  4288 => '0',
  4289 => '0',
  4290 => '0',
  4291 => '1',
  4292 => '1',
  4293 => '1',
  4294 => '1',
  4295 => '0',
  4296 => '0',
  4297 => '0',
  4298 => '1',
  4299 => '1',
  4300 => '0',
  4301 => '0',
  4302 => '0',
  4303 => '0',
  4304 => '0',
  4305 => '1',
  4306 => '1',
  4307 => '0',
  4308 => '0',
  4309 => '0',
  4310 => '0',
  4311 => '0',
  4312 => '0',
  4313 => '1',
  4314 => '1',
  4315 => '0',
  4316 => '0',
  4317 => '0',
  4318 => '0',
  4319 => '0',
  4320 => '0',
  4321 => '1',
  4322 => '1',
  4323 => '0',
  4324 => '0',
  4325 => '0',
  4326 => '0',
  4327 => '0',
  4328 => '0',
  4329 => '0',
  4330 => '1',
  4331 => '1',
  4332 => '0',
  4333 => '0',
  4334 => '0',
  4335 => '0',
  4336 => '0',
  4337 => '0',
  4338 => '0',
  4339 => '1',
  4340 => '1',
  4341 => '1',
  4342 => '1',
  4343 => '0',
  4344 => '0',
  4345 => '0',
  4346 => '0',
  4347 => '0',
  4348 => '0',
  4349 => '0',
  4350 => '0',
  4351 => '0',
  4352 => '0',
  4353 => '1',
  4354 => '1',
  4355 => '1',
  4356 => '1',
  4357 => '0',
  4358 => '0',
  4359 => '0',
  4360 => '0',
  4361 => '1',
  4362 => '1',
  4363 => '0',
  4364 => '1',
  4365 => '1',
  4366 => '0',
  4367 => '0',
  4368 => '0',
  4369 => '1',
  4370 => '1',
  4371 => '0',
  4372 => '0',
  4373 => '1',
  4374 => '1',
  4375 => '0',
  4376 => '0',
  4377 => '1',
  4378 => '1',
  4379 => '0',
  4380 => '0',
  4381 => '1',
  4382 => '1',
  4383 => '0',
  4384 => '0',
  4385 => '1',
  4386 => '1',
  4387 => '0',
  4388 => '0',
  4389 => '1',
  4390 => '1',
  4391 => '0',
  4392 => '0',
  4393 => '1',
  4394 => '1',
  4395 => '0',
  4396 => '1',
  4397 => '1',
  4398 => '0',
  4399 => '0',
  4400 => '0',
  4401 => '1',
  4402 => '1',
  4403 => '1',
  4404 => '1',
  4405 => '0',
  4406 => '0',
  4407 => '0',
  4408 => '0',
  4409 => '0',
  4410 => '0',
  4411 => '0',
  4412 => '0',
  4413 => '0',
  4414 => '0',
  4415 => '0',
  4416 => '0',
  4417 => '1',
  4418 => '1',
  4419 => '1',
  4420 => '1',
  4421 => '1',
  4422 => '1',
  4423 => '0',
  4424 => '0',
  4425 => '1',
  4426 => '1',
  4427 => '0',
  4428 => '0',
  4429 => '0',
  4430 => '0',
  4431 => '0',
  4432 => '0',
  4433 => '1',
  4434 => '1',
  4435 => '0',
  4436 => '0',
  4437 => '0',
  4438 => '0',
  4439 => '0',
  4440 => '0',
  4441 => '1',
  4442 => '1',
  4443 => '1',
  4444 => '1',
  4445 => '0',
  4446 => '0',
  4447 => '0',
  4448 => '0',
  4449 => '1',
  4450 => '1',
  4451 => '0',
  4452 => '0',
  4453 => '0',
  4454 => '0',
  4455 => '0',
  4456 => '0',
  4457 => '1',
  4458 => '1',
  4459 => '0',
  4460 => '0',
  4461 => '0',
  4462 => '0',
  4463 => '0',
  4464 => '0',
  4465 => '1',
  4466 => '1',
  4467 => '1',
  4468 => '1',
  4469 => '1',
  4470 => '1',
  4471 => '0',
  4472 => '0',
  4473 => '0',
  4474 => '0',
  4475 => '0',
  4476 => '0',
  4477 => '0',
  4478 => '0',
  4479 => '0',
  4480 => '0',
  4481 => '1',
  4482 => '1',
  4483 => '1',
  4484 => '1',
  4485 => '1',
  4486 => '1',
  4487 => '0',
  4488 => '0',
  4489 => '1',
  4490 => '1',
  4491 => '0',
  4492 => '0',
  4493 => '0',
  4494 => '0',
  4495 => '0',
  4496 => '0',
  4497 => '1',
  4498 => '1',
  4499 => '0',
  4500 => '0',
  4501 => '0',
  4502 => '0',
  4503 => '0',
  4504 => '0',
  4505 => '1',
  4506 => '1',
  4507 => '1',
  4508 => '1',
  4509 => '0',
  4510 => '0',
  4511 => '0',
  4512 => '0',
  4513 => '1',
  4514 => '1',
  4515 => '0',
  4516 => '0',
  4517 => '0',
  4518 => '0',
  4519 => '0',
  4520 => '0',
  4521 => '1',
  4522 => '1',
  4523 => '0',
  4524 => '0',
  4525 => '0',
  4526 => '0',
  4527 => '0',
  4528 => '0',
  4529 => '1',
  4530 => '1',
  4531 => '0',
  4532 => '0',
  4533 => '0',
  4534 => '0',
  4535 => '0',
  4536 => '0',
  4537 => '0',
  4538 => '0',
  4539 => '0',
  4540 => '0',
  4541 => '0',
  4542 => '0',
  4543 => '0',
  4544 => '0',
  4545 => '0',
  4546 => '1',
  4547 => '1',
  4548 => '1',
  4549 => '1',
  4550 => '0',
  4551 => '0',
  4552 => '0',
  4553 => '1',
  4554 => '1',
  4555 => '0',
  4556 => '0',
  4557 => '1',
  4558 => '1',
  4559 => '0',
  4560 => '0',
  4561 => '1',
  4562 => '1',
  4563 => '0',
  4564 => '0',
  4565 => '0',
  4566 => '0',
  4567 => '0',
  4568 => '0',
  4569 => '1',
  4570 => '1',
  4571 => '0',
  4572 => '1',
  4573 => '1',
  4574 => '1',
  4575 => '0',
  4576 => '0',
  4577 => '1',
  4578 => '1',
  4579 => '0',
  4580 => '0',
  4581 => '1',
  4582 => '1',
  4583 => '0',
  4584 => '0',
  4585 => '1',
  4586 => '1',
  4587 => '0',
  4588 => '0',
  4589 => '1',
  4590 => '1',
  4591 => '0',
  4592 => '0',
  4593 => '0',
  4594 => '1',
  4595 => '1',
  4596 => '1',
  4597 => '1',
  4598 => '1',
  4599 => '0',
  4600 => '0',
  4601 => '0',
  4602 => '0',
  4603 => '0',
  4604 => '0',
  4605 => '0',
  4606 => '0',
  4607 => '0',
  4608 => '0',
  4609 => '1',
  4610 => '1',
  4611 => '0',
  4612 => '0',
  4613 => '1',
  4614 => '1',
  4615 => '0',
  4616 => '0',
  4617 => '1',
  4618 => '1',
  4619 => '0',
  4620 => '0',
  4621 => '1',
  4622 => '1',
  4623 => '0',
  4624 => '0',
  4625 => '1',
  4626 => '1',
  4627 => '0',
  4628 => '0',
  4629 => '1',
  4630 => '1',
  4631 => '0',
  4632 => '0',
  4633 => '1',
  4634 => '1',
  4635 => '1',
  4636 => '1',
  4637 => '1',
  4638 => '1',
  4639 => '0',
  4640 => '0',
  4641 => '1',
  4642 => '1',
  4643 => '0',
  4644 => '0',
  4645 => '1',
  4646 => '1',
  4647 => '0',
  4648 => '0',
  4649 => '1',
  4650 => '1',
  4651 => '0',
  4652 => '0',
  4653 => '1',
  4654 => '1',
  4655 => '0',
  4656 => '0',
  4657 => '1',
  4658 => '1',
  4659 => '0',
  4660 => '0',
  4661 => '1',
  4662 => '1',
  4663 => '0',
  4664 => '0',
  4665 => '0',
  4666 => '0',
  4667 => '0',
  4668 => '0',
  4669 => '0',
  4670 => '0',
  4671 => '0',
  4672 => '0',
  4673 => '0',
  4674 => '1',
  4675 => '1',
  4676 => '1',
  4677 => '1',
  4678 => '0',
  4679 => '0',
  4680 => '0',
  4681 => '0',
  4682 => '0',
  4683 => '1',
  4684 => '1',
  4685 => '0',
  4686 => '0',
  4687 => '0',
  4688 => '0',
  4689 => '0',
  4690 => '0',
  4691 => '1',
  4692 => '1',
  4693 => '0',
  4694 => '0',
  4695 => '0',
  4696 => '0',
  4697 => '0',
  4698 => '0',
  4699 => '1',
  4700 => '1',
  4701 => '0',
  4702 => '0',
  4703 => '0',
  4704 => '0',
  4705 => '0',
  4706 => '0',
  4707 => '1',
  4708 => '1',
  4709 => '0',
  4710 => '0',
  4711 => '0',
  4712 => '0',
  4713 => '0',
  4714 => '0',
  4715 => '1',
  4716 => '1',
  4717 => '0',
  4718 => '0',
  4719 => '0',
  4720 => '0',
  4721 => '0',
  4722 => '1',
  4723 => '1',
  4724 => '1',
  4725 => '1',
  4726 => '0',
  4727 => '0',
  4728 => '0',
  4729 => '0',
  4730 => '0',
  4731 => '0',
  4732 => '0',
  4733 => '0',
  4734 => '0',
  4735 => '0',
  4736 => '0',
  4737 => '0',
  4738 => '0',
  4739 => '0',
  4740 => '0',
  4741 => '1',
  4742 => '1',
  4743 => '0',
  4744 => '0',
  4745 => '0',
  4746 => '0',
  4747 => '0',
  4748 => '0',
  4749 => '1',
  4750 => '1',
  4751 => '0',
  4752 => '0',
  4753 => '0',
  4754 => '0',
  4755 => '0',
  4756 => '0',
  4757 => '1',
  4758 => '1',
  4759 => '0',
  4760 => '0',
  4761 => '0',
  4762 => '0',
  4763 => '0',
  4764 => '0',
  4765 => '1',
  4766 => '1',
  4767 => '0',
  4768 => '0',
  4769 => '0',
  4770 => '0',
  4771 => '0',
  4772 => '0',
  4773 => '1',
  4774 => '1',
  4775 => '0',
  4776 => '0',
  4777 => '1',
  4778 => '1',
  4779 => '0',
  4780 => '0',
  4781 => '1',
  4782 => '1',
  4783 => '0',
  4784 => '0',
  4785 => '0',
  4786 => '1',
  4787 => '1',
  4788 => '1',
  4789 => '1',
  4790 => '0',
  4791 => '0',
  4792 => '0',
  4793 => '0',
  4794 => '0',
  4795 => '0',
  4796 => '0',
  4797 => '0',
  4798 => '0',
  4799 => '0',
  4800 => '1',
  4801 => '1',
  4802 => '0',
  4803 => '0',
  4804 => '0',
  4805 => '1',
  4806 => '1',
  4807 => '0',
  4808 => '1',
  4809 => '1',
  4810 => '0',
  4811 => '0',
  4812 => '1',
  4813 => '1',
  4814 => '0',
  4815 => '0',
  4816 => '1',
  4817 => '1',
  4818 => '0',
  4819 => '1',
  4820 => '1',
  4821 => '0',
  4822 => '0',
  4823 => '0',
  4824 => '1',
  4825 => '1',
  4826 => '1',
  4827 => '1',
  4828 => '0',
  4829 => '0',
  4830 => '0',
  4831 => '0',
  4832 => '1',
  4833 => '1',
  4834 => '0',
  4835 => '1',
  4836 => '1',
  4837 => '0',
  4838 => '0',
  4839 => '0',
  4840 => '1',
  4841 => '1',
  4842 => '0',
  4843 => '0',
  4844 => '1',
  4845 => '1',
  4846 => '0',
  4847 => '0',
  4848 => '1',
  4849 => '1',
  4850 => '0',
  4851 => '0',
  4852 => '0',
  4853 => '1',
  4854 => '1',
  4855 => '0',
  4856 => '0',
  4857 => '0',
  4858 => '0',
  4859 => '0',
  4860 => '0',
  4861 => '0',
  4862 => '0',
  4863 => '0',
  4864 => '0',
  4865 => '1',
  4866 => '1',
  4867 => '0',
  4868 => '0',
  4869 => '0',
  4870 => '0',
  4871 => '0',
  4872 => '0',
  4873 => '1',
  4874 => '1',
  4875 => '0',
  4876 => '0',
  4877 => '0',
  4878 => '0',
  4879 => '0',
  4880 => '0',
  4881 => '1',
  4882 => '1',
  4883 => '0',
  4884 => '0',
  4885 => '0',
  4886 => '0',
  4887 => '0',
  4888 => '0',
  4889 => '1',
  4890 => '1',
  4891 => '0',
  4892 => '0',
  4893 => '0',
  4894 => '0',
  4895 => '0',
  4896 => '0',
  4897 => '1',
  4898 => '1',
  4899 => '0',
  4900 => '0',
  4901 => '0',
  4902 => '0',
  4903 => '0',
  4904 => '0',
  4905 => '1',
  4906 => '1',
  4907 => '0',
  4908 => '0',
  4909 => '0',
  4910 => '0',
  4911 => '0',
  4912 => '0',
  4913 => '1',
  4914 => '1',
  4915 => '1',
  4916 => '1',
  4917 => '1',
  4918 => '1',
  4919 => '0',
  4920 => '0',
  4921 => '0',
  4922 => '0',
  4923 => '0',
  4924 => '0',
  4925 => '0',
  4926 => '0',
  4927 => '0',
  4928 => '1',
  4929 => '1',
  4930 => '0',
  4931 => '0',
  4932 => '0',
  4933 => '1',
  4934 => '1',
  4935 => '0',
  4936 => '1',
  4937 => '1',
  4938 => '1',
  4939 => '0',
  4940 => '1',
  4941 => '1',
  4942 => '1',
  4943 => '0',
  4944 => '1',
  4945 => '1',
  4946 => '1',
  4947 => '1',
  4948 => '1',
  4949 => '1',
  4950 => '1',
  4951 => '0',
  4952 => '1',
  4953 => '1',
  4954 => '0',
  4955 => '1',
  4956 => '0',
  4957 => '1',
  4958 => '1',
  4959 => '0',
  4960 => '1',
  4961 => '1',
  4962 => '0',
  4963 => '0',
  4964 => '0',
  4965 => '1',
  4966 => '1',
  4967 => '0',
  4968 => '1',
  4969 => '1',
  4970 => '0',
  4971 => '0',
  4972 => '0',
  4973 => '1',
  4974 => '1',
  4975 => '0',
  4976 => '1',
  4977 => '1',
  4978 => '0',
  4979 => '0',
  4980 => '0',
  4981 => '1',
  4982 => '1',
  4983 => '0',
  4984 => '0',
  4985 => '0',
  4986 => '0',
  4987 => '0',
  4988 => '0',
  4989 => '0',
  4990 => '0',
  4991 => '0',
  4992 => '1',
  4993 => '1',
  4994 => '0',
  4995 => '0',
  4996 => '0',
  4997 => '1',
  4998 => '1',
  4999 => '0',
  5000 => '1',
  5001 => '1',
  5002 => '1',
  5003 => '0',
  5004 => '0',
  5005 => '1',
  5006 => '1',
  5007 => '0',
  5008 => '1',
  5009 => '1',
  5010 => '1',
  5011 => '1',
  5012 => '0',
  5013 => '1',
  5014 => '1',
  5015 => '0',
  5016 => '1',
  5017 => '1',
  5018 => '0',
  5019 => '1',
  5020 => '1',
  5021 => '1',
  5022 => '1',
  5023 => '0',
  5024 => '1',
  5025 => '1',
  5026 => '0',
  5027 => '0',
  5028 => '1',
  5029 => '1',
  5030 => '1',
  5031 => '0',
  5032 => '1',
  5033 => '1',
  5034 => '0',
  5035 => '0',
  5036 => '0',
  5037 => '1',
  5038 => '1',
  5039 => '0',
  5040 => '1',
  5041 => '1',
  5042 => '0',
  5043 => '0',
  5044 => '0',
  5045 => '1',
  5046 => '1',
  5047 => '0',
  5048 => '0',
  5049 => '0',
  5050 => '0',
  5051 => '0',
  5052 => '0',
  5053 => '0',
  5054 => '0',
  5055 => '0',
  5056 => '0',
  5057 => '0',
  5058 => '1',
  5059 => '1',
  5060 => '1',
  5061 => '1',
  5062 => '0',
  5063 => '0',
  5064 => '0',
  5065 => '1',
  5066 => '1',
  5067 => '0',
  5068 => '0',
  5069 => '1',
  5070 => '1',
  5071 => '0',
  5072 => '0',
  5073 => '1',
  5074 => '1',
  5075 => '0',
  5076 => '0',
  5077 => '1',
  5078 => '1',
  5079 => '0',
  5080 => '0',
  5081 => '1',
  5082 => '1',
  5083 => '0',
  5084 => '0',
  5085 => '1',
  5086 => '1',
  5087 => '0',
  5088 => '0',
  5089 => '1',
  5090 => '1',
  5091 => '0',
  5092 => '0',
  5093 => '1',
  5094 => '1',
  5095 => '0',
  5096 => '0',
  5097 => '1',
  5098 => '1',
  5099 => '0',
  5100 => '0',
  5101 => '1',
  5102 => '1',
  5103 => '0',
  5104 => '0',
  5105 => '0',
  5106 => '1',
  5107 => '1',
  5108 => '1',
  5109 => '1',
  5110 => '0',
  5111 => '0',
  5112 => '0',
  5113 => '0',
  5114 => '0',
  5115 => '0',
  5116 => '0',
  5117 => '0',
  5118 => '0',
  5119 => '0',
  5120 => '0',
  5121 => '1',
  5122 => '1',
  5123 => '1',
  5124 => '1',
  5125 => '1',
  5126 => '0',
  5127 => '0',
  5128 => '0',
  5129 => '1',
  5130 => '1',
  5131 => '0',
  5132 => '0',
  5133 => '1',
  5134 => '1',
  5135 => '0',
  5136 => '0',
  5137 => '1',
  5138 => '1',
  5139 => '0',
  5140 => '0',
  5141 => '1',
  5142 => '1',
  5143 => '0',
  5144 => '0',
  5145 => '1',
  5146 => '1',
  5147 => '1',
  5148 => '1',
  5149 => '1',
  5150 => '0',
  5151 => '0',
  5152 => '0',
  5153 => '1',
  5154 => '1',
  5155 => '0',
  5156 => '0',
  5157 => '0',
  5158 => '0',
  5159 => '0',
  5160 => '0',
  5161 => '1',
  5162 => '1',
  5163 => '0',
  5164 => '0',
  5165 => '0',
  5166 => '0',
  5167 => '0',
  5168 => '0',
  5169 => '1',
  5170 => '1',
  5171 => '0',
  5172 => '0',
  5173 => '0',
  5174 => '0',
  5175 => '0',
  5176 => '0',
  5177 => '0',
  5178 => '0',
  5179 => '0',
  5180 => '0',
  5181 => '0',
  5182 => '0',
  5183 => '0',
  5184 => '0',
  5185 => '1',
  5186 => '1',
  5187 => '1',
  5188 => '1',
  5189 => '0',
  5190 => '0',
  5191 => '0',
  5192 => '1',
  5193 => '1',
  5194 => '0',
  5195 => '0',
  5196 => '1',
  5197 => '1',
  5198 => '0',
  5199 => '0',
  5200 => '1',
  5201 => '1',
  5202 => '0',
  5203 => '0',
  5204 => '1',
  5205 => '1',
  5206 => '0',
  5207 => '0',
  5208 => '1',
  5209 => '1',
  5210 => '0',
  5211 => '0',
  5212 => '1',
  5213 => '1',
  5214 => '0',
  5215 => '0',
  5216 => '1',
  5217 => '1',
  5218 => '0',
  5219 => '0',
  5220 => '1',
  5221 => '1',
  5222 => '0',
  5223 => '0',
  5224 => '1',
  5225 => '1',
  5226 => '0',
  5227 => '1',
  5228 => '1',
  5229 => '1',
  5230 => '0',
  5231 => '0',
  5232 => '0',
  5233 => '1',
  5234 => '1',
  5235 => '1',
  5236 => '1',
  5237 => '1',
  5238 => '1',
  5239 => '0',
  5240 => '0',
  5241 => '0',
  5242 => '0',
  5243 => '0',
  5244 => '0',
  5245 => '0',
  5246 => '0',
  5247 => '0',
  5248 => '0',
  5249 => '1',
  5250 => '1',
  5251 => '1',
  5252 => '1',
  5253 => '1',
  5254 => '0',
  5255 => '0',
  5256 => '0',
  5257 => '1',
  5258 => '1',
  5259 => '0',
  5260 => '0',
  5261 => '1',
  5262 => '1',
  5263 => '0',
  5264 => '0',
  5265 => '1',
  5266 => '1',
  5267 => '0',
  5268 => '0',
  5269 => '1',
  5270 => '1',
  5271 => '0',
  5272 => '0',
  5273 => '1',
  5274 => '1',
  5275 => '1',
  5276 => '1',
  5277 => '1',
  5278 => '0',
  5279 => '0',
  5280 => '0',
  5281 => '1',
  5282 => '1',
  5283 => '0',
  5284 => '1',
  5285 => '1',
  5286 => '0',
  5287 => '0',
  5288 => '0',
  5289 => '1',
  5290 => '1',
  5291 => '0',
  5292 => '0',
  5293 => '1',
  5294 => '1',
  5295 => '0',
  5296 => '0',
  5297 => '1',
  5298 => '1',
  5299 => '0',
  5300 => '0',
  5301 => '1',
  5302 => '1',
  5303 => '0',
  5304 => '0',
  5305 => '0',
  5306 => '0',
  5307 => '0',
  5308 => '0',
  5309 => '0',
  5310 => '0',
  5311 => '0',
  5312 => '0',
  5313 => '0',
  5314 => '1',
  5315 => '1',
  5316 => '1',
  5317 => '1',
  5318 => '0',
  5319 => '0',
  5320 => '0',
  5321 => '1',
  5322 => '1',
  5323 => '0',
  5324 => '0',
  5325 => '1',
  5326 => '1',
  5327 => '0',
  5328 => '0',
  5329 => '1',
  5330 => '1',
  5331 => '1',
  5332 => '0',
  5333 => '0',
  5334 => '0',
  5335 => '0',
  5336 => '0',
  5337 => '0',
  5338 => '1',
  5339 => '1',
  5340 => '1',
  5341 => '1',
  5342 => '0',
  5343 => '0',
  5344 => '0',
  5345 => '0',
  5346 => '0',
  5347 => '0',
  5348 => '1',
  5349 => '1',
  5350 => '1',
  5351 => '0',
  5352 => '0',
  5353 => '1',
  5354 => '1',
  5355 => '0',
  5356 => '0',
  5357 => '1',
  5358 => '1',
  5359 => '0',
  5360 => '0',
  5361 => '0',
  5362 => '1',
  5363 => '1',
  5364 => '1',
  5365 => '1',
  5366 => '0',
  5367 => '0',
  5368 => '0',
  5369 => '0',
  5370 => '0',
  5371 => '0',
  5372 => '0',
  5373 => '0',
  5374 => '0',
  5375 => '0',
  5376 => '0',
  5377 => '1',
  5378 => '1',
  5379 => '1',
  5380 => '1',
  5381 => '1',
  5382 => '1',
  5383 => '0',
  5384 => '0',
  5385 => '0',
  5386 => '0',
  5387 => '1',
  5388 => '1',
  5389 => '0',
  5390 => '0',
  5391 => '0',
  5392 => '0',
  5393 => '0',
  5394 => '0',
  5395 => '1',
  5396 => '1',
  5397 => '0',
  5398 => '0',
  5399 => '0',
  5400 => '0',
  5401 => '0',
  5402 => '0',
  5403 => '1',
  5404 => '1',
  5405 => '0',
  5406 => '0',
  5407 => '0',
  5408 => '0',
  5409 => '0',
  5410 => '0',
  5411 => '1',
  5412 => '1',
  5413 => '0',
  5414 => '0',
  5415 => '0',
  5416 => '0',
  5417 => '0',
  5418 => '0',
  5419 => '1',
  5420 => '1',
  5421 => '0',
  5422 => '0',
  5423 => '0',
  5424 => '0',
  5425 => '0',
  5426 => '0',
  5427 => '1',
  5428 => '1',
  5429 => '0',
  5430 => '0',
  5431 => '0',
  5432 => '0',
  5433 => '0',
  5434 => '0',
  5435 => '0',
  5436 => '0',
  5437 => '0',
  5438 => '0',
  5439 => '0',
  5440 => '0',
  5441 => '1',
  5442 => '1',
  5443 => '0',
  5444 => '0',
  5445 => '1',
  5446 => '1',
  5447 => '0',
  5448 => '0',
  5449 => '1',
  5450 => '1',
  5451 => '0',
  5452 => '0',
  5453 => '1',
  5454 => '1',
  5455 => '0',
  5456 => '0',
  5457 => '1',
  5458 => '1',
  5459 => '0',
  5460 => '0',
  5461 => '1',
  5462 => '1',
  5463 => '0',
  5464 => '0',
  5465 => '1',
  5466 => '1',
  5467 => '0',
  5468 => '0',
  5469 => '1',
  5470 => '1',
  5471 => '0',
  5472 => '0',
  5473 => '1',
  5474 => '1',
  5475 => '0',
  5476 => '0',
  5477 => '1',
  5478 => '1',
  5479 => '0',
  5480 => '0',
  5481 => '1',
  5482 => '1',
  5483 => '0',
  5484 => '0',
  5485 => '1',
  5486 => '1',
  5487 => '0',
  5488 => '0',
  5489 => '0',
  5490 => '1',
  5491 => '1',
  5492 => '1',
  5493 => '1',
  5494 => '0',
  5495 => '0',
  5496 => '0',
  5497 => '0',
  5498 => '0',
  5499 => '0',
  5500 => '0',
  5501 => '0',
  5502 => '0',
  5503 => '0',
  5504 => '0',
  5505 => '1',
  5506 => '1',
  5507 => '0',
  5508 => '0',
  5509 => '1',
  5510 => '1',
  5511 => '0',
  5512 => '0',
  5513 => '1',
  5514 => '1',
  5515 => '0',
  5516 => '0',
  5517 => '1',
  5518 => '1',
  5519 => '0',
  5520 => '0',
  5521 => '1',
  5522 => '1',
  5523 => '0',
  5524 => '0',
  5525 => '1',
  5526 => '1',
  5527 => '0',
  5528 => '0',
  5529 => '1',
  5530 => '1',
  5531 => '0',
  5532 => '0',
  5533 => '1',
  5534 => '1',
  5535 => '0',
  5536 => '0',
  5537 => '0',
  5538 => '1',
  5539 => '1',
  5540 => '1',
  5541 => '1',
  5542 => '0',
  5543 => '0',
  5544 => '0',
  5545 => '0',
  5546 => '1',
  5547 => '1',
  5548 => '1',
  5549 => '1',
  5550 => '0',
  5551 => '0',
  5552 => '0',
  5553 => '0',
  5554 => '0',
  5555 => '1',
  5556 => '1',
  5557 => '0',
  5558 => '0',
  5559 => '0',
  5560 => '0',
  5561 => '0',
  5562 => '0',
  5563 => '0',
  5564 => '0',
  5565 => '0',
  5566 => '0',
  5567 => '0',
  5568 => '1',
  5569 => '1',
  5570 => '0',
  5571 => '0',
  5572 => '0',
  5573 => '1',
  5574 => '1',
  5575 => '0',
  5576 => '1',
  5577 => '1',
  5578 => '0',
  5579 => '0',
  5580 => '0',
  5581 => '1',
  5582 => '1',
  5583 => '0',
  5584 => '1',
  5585 => '1',
  5586 => '0',
  5587 => '0',
  5588 => '0',
  5589 => '1',
  5590 => '1',
  5591 => '0',
  5592 => '1',
  5593 => '1',
  5594 => '0',
  5595 => '1',
  5596 => '0',
  5597 => '1',
  5598 => '1',
  5599 => '0',
  5600 => '1',
  5601 => '1',
  5602 => '1',
  5603 => '1',
  5604 => '1',
  5605 => '1',
  5606 => '1',
  5607 => '0',
  5608 => '1',
  5609 => '1',
  5610 => '1',
  5611 => '0',
  5612 => '1',
  5613 => '1',
  5614 => '1',
  5615 => '0',
  5616 => '1',
  5617 => '1',
  5618 => '0',
  5619 => '0',
  5620 => '0',
  5621 => '1',
  5622 => '1',
  5623 => '0',
  5624 => '0',
  5625 => '0',
  5626 => '0',
  5627 => '0',
  5628 => '0',
  5629 => '0',
  5630 => '0',
  5631 => '0',
  5632 => '1',
  5633 => '1',
  5634 => '0',
  5635 => '0',
  5636 => '0',
  5637 => '0',
  5638 => '1',
  5639 => '1',
  5640 => '0',
  5641 => '1',
  5642 => '1',
  5643 => '0',
  5644 => '0',
  5645 => '1',
  5646 => '1',
  5647 => '0',
  5648 => '0',
  5649 => '0',
  5650 => '1',
  5651 => '1',
  5652 => '1',
  5653 => '1',
  5654 => '0',
  5655 => '0',
  5656 => '0',
  5657 => '0',
  5658 => '0',
  5659 => '1',
  5660 => '1',
  5661 => '0',
  5662 => '0',
  5663 => '0',
  5664 => '0',
  5665 => '0',
  5666 => '1',
  5667 => '1',
  5668 => '1',
  5669 => '1',
  5670 => '0',
  5671 => '0',
  5672 => '0',
  5673 => '1',
  5674 => '1',
  5675 => '0',
  5676 => '0',
  5677 => '1',
  5678 => '1',
  5679 => '0',
  5680 => '1',
  5681 => '1',
  5682 => '0',
  5683 => '0',
  5684 => '0',
  5685 => '0',
  5686 => '1',
  5687 => '1',
  5688 => '0',
  5689 => '0',
  5690 => '0',
  5691 => '0',
  5692 => '0',
  5693 => '0',
  5694 => '0',
  5695 => '0',
  5696 => '1',
  5697 => '1',
  5698 => '0',
  5699 => '0',
  5700 => '0',
  5701 => '0',
  5702 => '1',
  5703 => '1',
  5704 => '0',
  5705 => '1',
  5706 => '1',
  5707 => '0',
  5708 => '0',
  5709 => '1',
  5710 => '1',
  5711 => '0',
  5712 => '0',
  5713 => '0',
  5714 => '1',
  5715 => '1',
  5716 => '1',
  5717 => '1',
  5718 => '0',
  5719 => '0',
  5720 => '0',
  5721 => '0',
  5722 => '0',
  5723 => '1',
  5724 => '1',
  5725 => '0',
  5726 => '0',
  5727 => '0',
  5728 => '0',
  5729 => '0',
  5730 => '0',
  5731 => '1',
  5732 => '1',
  5733 => '0',
  5734 => '0',
  5735 => '0',
  5736 => '0',
  5737 => '0',
  5738 => '0',
  5739 => '1',
  5740 => '1',
  5741 => '0',
  5742 => '0',
  5743 => '0',
  5744 => '0',
  5745 => '0',
  5746 => '0',
  5747 => '1',
  5748 => '1',
  5749 => '0',
  5750 => '0',
  5751 => '0',
  5752 => '0',
  5753 => '0',
  5754 => '0',
  5755 => '0',
  5756 => '0',
  5757 => '0',
  5758 => '0',
  5759 => '0',
  5760 => '1',
  5761 => '1',
  5762 => '1',
  5763 => '1',
  5764 => '1',
  5765 => '1',
  5766 => '1',
  5767 => '0',
  5768 => '0',
  5769 => '0',
  5770 => '0',
  5771 => '0',
  5772 => '1',
  5773 => '1',
  5774 => '0',
  5775 => '0',
  5776 => '0',
  5777 => '0',
  5778 => '0',
  5779 => '1',
  5780 => '1',
  5781 => '0',
  5782 => '0',
  5783 => '0',
  5784 => '0',
  5785 => '0',
  5786 => '1',
  5787 => '1',
  5788 => '0',
  5789 => '0',
  5790 => '0',
  5791 => '0',
  5792 => '0',
  5793 => '1',
  5794 => '1',
  5795 => '0',
  5796 => '0',
  5797 => '0',
  5798 => '0',
  5799 => '0',
  5800 => '1',
  5801 => '1',
  5802 => '0',
  5803 => '0',
  5804 => '0',
  5805 => '0',
  5806 => '0',
  5807 => '0',
  5808 => '1',
  5809 => '1',
  5810 => '1',
  5811 => '1',
  5812 => '1',
  5813 => '1',
  5814 => '1',
  5815 => '0',
  5816 => '0',
  5817 => '0',
  5818 => '0',
  5819 => '0',
  5820 => '0',
  5821 => '0',
  5822 => '0',
  5823 => '0',
  5824 => '0',
  5825 => '0',
  5826 => '1',
  5827 => '1',
  5828 => '1',
  5829 => '1',
  5830 => '0',
  5831 => '0',
  5832 => '0',
  5833 => '0',
  5834 => '1',
  5835 => '1',
  5836 => '0',
  5837 => '0',
  5838 => '0',
  5839 => '0',
  5840 => '0',
  5841 => '0',
  5842 => '1',
  5843 => '1',
  5844 => '0',
  5845 => '0',
  5846 => '0',
  5847 => '0',
  5848 => '0',
  5849 => '0',
  5850 => '1',
  5851 => '1',
  5852 => '0',
  5853 => '0',
  5854 => '0',
  5855 => '0',
  5856 => '0',
  5857 => '0',
  5858 => '1',
  5859 => '1',
  5860 => '0',
  5861 => '0',
  5862 => '0',
  5863 => '0',
  5864 => '0',
  5865 => '0',
  5866 => '1',
  5867 => '1',
  5868 => '0',
  5869 => '0',
  5870 => '0',
  5871 => '0',
  5872 => '0',
  5873 => '0',
  5874 => '1',
  5875 => '1',
  5876 => '1',
  5877 => '1',
  5878 => '0',
  5879 => '0',
  5880 => '0',
  5881 => '0',
  5882 => '0',
  5883 => '0',
  5884 => '0',
  5885 => '0',
  5886 => '0',
  5887 => '0',
  5888 => '1',
  5889 => '1',
  5890 => '0',
  5891 => '0',
  5892 => '0',
  5893 => '0',
  5894 => '0',
  5895 => '0',
  5896 => '0',
  5897 => '1',
  5898 => '1',
  5899 => '0',
  5900 => '0',
  5901 => '0',
  5902 => '0',
  5903 => '0',
  5904 => '0',
  5905 => '0',
  5906 => '1',
  5907 => '1',
  5908 => '0',
  5909 => '0',
  5910 => '0',
  5911 => '0',
  5912 => '0',
  5913 => '0',
  5914 => '0',
  5915 => '1',
  5916 => '1',
  5917 => '0',
  5918 => '0',
  5919 => '0',
  5920 => '0',
  5921 => '0',
  5922 => '0',
  5923 => '0',
  5924 => '1',
  5925 => '1',
  5926 => '0',
  5927 => '0',
  5928 => '0',
  5929 => '0',
  5930 => '0',
  5931 => '0',
  5932 => '0',
  5933 => '1',
  5934 => '1',
  5935 => '0',
  5936 => '0',
  5937 => '0',
  5938 => '0',
  5939 => '0',
  5940 => '0',
  5941 => '0',
  5942 => '1',
  5943 => '1',
  5944 => '0',
  5945 => '0',
  5946 => '0',
  5947 => '0',
  5948 => '0',
  5949 => '0',
  5950 => '0',
  5951 => '0',
  5952 => '0',
  5953 => '0',
  5954 => '1',
  5955 => '1',
  5956 => '1',
  5957 => '1',
  5958 => '0',
  5959 => '0',
  5960 => '0',
  5961 => '0',
  5962 => '0',
  5963 => '0',
  5964 => '1',
  5965 => '1',
  5966 => '0',
  5967 => '0',
  5968 => '0',
  5969 => '0',
  5970 => '0',
  5971 => '0',
  5972 => '1',
  5973 => '1',
  5974 => '0',
  5975 => '0',
  5976 => '0',
  5977 => '0',
  5978 => '0',
  5979 => '0',
  5980 => '1',
  5981 => '1',
  5982 => '0',
  5983 => '0',
  5984 => '0',
  5985 => '0',
  5986 => '0',
  5987 => '0',
  5988 => '1',
  5989 => '1',
  5990 => '0',
  5991 => '0',
  5992 => '0',
  5993 => '0',
  5994 => '0',
  5995 => '0',
  5996 => '1',
  5997 => '1',
  5998 => '0',
  5999 => '0',
  6000 => '0',
  6001 => '0',
  6002 => '1',
  6003 => '1',
  6004 => '1',
  6005 => '1',
  6006 => '0',
  6007 => '0',
  6008 => '0',
  6009 => '0',
  6010 => '0',
  6011 => '0',
  6012 => '0',
  6013 => '0',
  6014 => '0',
  6015 => '0',
  6016 => '0',
  6017 => '0',
  6018 => '0',
  6019 => '1',
  6020 => '0',
  6021 => '0',
  6022 => '0',
  6023 => '0',
  6024 => '0',
  6025 => '0',
  6026 => '1',
  6027 => '1',
  6028 => '1',
  6029 => '0',
  6030 => '0',
  6031 => '0',
  6032 => '0',
  6033 => '1',
  6034 => '1',
  6035 => '0',
  6036 => '1',
  6037 => '1',
  6038 => '0',
  6039 => '0',
  6040 => '1',
  6041 => '1',
  6042 => '0',
  6043 => '0',
  6044 => '0',
  6045 => '1',
  6046 => '1',
  6047 => '0',
  6048 => '0',
  6049 => '0',
  6050 => '0',
  6051 => '0',
  6052 => '0',
  6053 => '0',
  6054 => '0',
  6055 => '0',
  6056 => '0',
  6057 => '0',
  6058 => '0',
  6059 => '0',
  6060 => '0',
  6061 => '0',
  6062 => '0',
  6063 => '0',
  6064 => '0',
  6065 => '0',
  6066 => '0',
  6067 => '0',
  6068 => '0',
  6069 => '0',
  6070 => '0',
  6071 => '0',
  6072 => '0',
  6073 => '0',
  6074 => '0',
  6075 => '0',
  6076 => '0',
  6077 => '0',
  6078 => '0',
  6079 => '0',
  6080 => '0',
  6081 => '0',
  6082 => '0',
  6083 => '0',
  6084 => '0',
  6085 => '0',
  6086 => '0',
  6087 => '0',
  6088 => '0',
  6089 => '0',
  6090 => '0',
  6091 => '0',
  6092 => '0',
  6093 => '0',
  6094 => '0',
  6095 => '0',
  6096 => '0',
  6097 => '0',
  6098 => '0',
  6099 => '0',
  6100 => '0',
  6101 => '0',
  6102 => '0',
  6103 => '0',
  6104 => '0',
  6105 => '0',
  6106 => '0',
  6107 => '0',
  6108 => '0',
  6109 => '0',
  6110 => '0',
  6111 => '0',
  6112 => '0',
  6113 => '0',
  6114 => '0',
  6115 => '0',
  6116 => '0',
  6117 => '0',
  6118 => '0',
  6119 => '0',
  6120 => '0',
  6121 => '0',
  6122 => '0',
  6123 => '0',
  6124 => '0',
  6125 => '0',
  6126 => '0',
  6127 => '0',
  6128 => '0',
  6129 => '0',
  6130 => '0',
  6131 => '0',
  6132 => '0',
  6133 => '0',
  6134 => '0',
  6135 => '0',
  6136 => '1',
  6137 => '1',
  6138 => '1',
  6139 => '1',
  6140 => '1',
  6141 => '1',
  6142 => '1',
  6143 => '0',
  6144 => '0',
  6145 => '0',
  6146 => '0',
  6147 => '1',
  6148 => '1',
  6149 => '0',
  6150 => '0',
  6151 => '0',
  6152 => '0',
  6153 => '0',
  6154 => '0',
  6155 => '1',
  6156 => '1',
  6157 => '0',
  6158 => '0',
  6159 => '0',
  6160 => '0',
  6161 => '0',
  6162 => '0',
  6163 => '0',
  6164 => '1',
  6165 => '1',
  6166 => '0',
  6167 => '0',
  6168 => '0',
  6169 => '0',
  6170 => '0',
  6171 => '0',
  6172 => '0',
  6173 => '0',
  6174 => '0',
  6175 => '0',
  6176 => '0',
  6177 => '0',
  6178 => '0',
  6179 => '0',
  6180 => '0',
  6181 => '0',
  6182 => '0',
  6183 => '0',
  6184 => '0',
  6185 => '0',
  6186 => '0',
  6187 => '0',
  6188 => '0',
  6189 => '0',
  6190 => '0',
  6191 => '0',
  6192 => '0',
  6193 => '0',
  6194 => '0',
  6195 => '0',
  6196 => '0',
  6197 => '0',
  6198 => '0',
  6199 => '0',
  6200 => '0',
  6201 => '0',
  6202 => '0',
  6203 => '0',
  6204 => '0',
  6205 => '0',
  6206 => '0',
  6207 => '0',
  6208 => '0',
  6209 => '0',
  6210 => '0',
  6211 => '0',
  6212 => '0',
  6213 => '0',
  6214 => '0',
  6215 => '0',
  6216 => '0',
  6217 => '0',
  6218 => '0',
  6219 => '0',
  6220 => '0',
  6221 => '0',
  6222 => '0',
  6223 => '0',
  6224 => '0',
  6225 => '0',
  6226 => '1',
  6227 => '1',
  6228 => '1',
  6229 => '1',
  6230 => '0',
  6231 => '0',
  6232 => '0',
  6233 => '0',
  6234 => '0',
  6235 => '0',
  6236 => '0',
  6237 => '1',
  6238 => '1',
  6239 => '0',
  6240 => '0',
  6241 => '0',
  6242 => '1',
  6243 => '1',
  6244 => '1',
  6245 => '1',
  6246 => '1',
  6247 => '0',
  6248 => '0',
  6249 => '1',
  6250 => '1',
  6251 => '0',
  6252 => '0',
  6253 => '1',
  6254 => '1',
  6255 => '0',
  6256 => '0',
  6257 => '0',
  6258 => '1',
  6259 => '1',
  6260 => '1',
  6261 => '1',
  6262 => '1',
  6263 => '0',
  6264 => '0',
  6265 => '0',
  6266 => '0',
  6267 => '0',
  6268 => '0',
  6269 => '0',
  6270 => '0',
  6271 => '0',
  6272 => '0',
  6273 => '1',
  6274 => '1',
  6275 => '0',
  6276 => '0',
  6277 => '0',
  6278 => '0',
  6279 => '0',
  6280 => '0',
  6281 => '1',
  6282 => '1',
  6283 => '0',
  6284 => '0',
  6285 => '0',
  6286 => '0',
  6287 => '0',
  6288 => '0',
  6289 => '1',
  6290 => '1',
  6291 => '1',
  6292 => '1',
  6293 => '1',
  6294 => '0',
  6295 => '0',
  6296 => '0',
  6297 => '1',
  6298 => '1',
  6299 => '0',
  6300 => '0',
  6301 => '1',
  6302 => '1',
  6303 => '0',
  6304 => '0',
  6305 => '1',
  6306 => '1',
  6307 => '0',
  6308 => '0',
  6309 => '1',
  6310 => '1',
  6311 => '0',
  6312 => '0',
  6313 => '1',
  6314 => '1',
  6315 => '0',
  6316 => '0',
  6317 => '1',
  6318 => '1',
  6319 => '0',
  6320 => '0',
  6321 => '1',
  6322 => '1',
  6323 => '1',
  6324 => '1',
  6325 => '1',
  6326 => '0',
  6327 => '0',
  6328 => '0',
  6329 => '0',
  6330 => '0',
  6331 => '0',
  6332 => '0',
  6333 => '0',
  6334 => '0',
  6335 => '0',
  6336 => '0',
  6337 => '0',
  6338 => '0',
  6339 => '0',
  6340 => '0',
  6341 => '0',
  6342 => '0',
  6343 => '0',
  6344 => '0',
  6345 => '0',
  6346 => '0',
  6347 => '0',
  6348 => '0',
  6349 => '0',
  6350 => '0',
  6351 => '0',
  6352 => '0',
  6353 => '0',
  6354 => '1',
  6355 => '1',
  6356 => '1',
  6357 => '1',
  6358 => '0',
  6359 => '0',
  6360 => '0',
  6361 => '1',
  6362 => '1',
  6363 => '0',
  6364 => '0',
  6365 => '0',
  6366 => '0',
  6367 => '0',
  6368 => '0',
  6369 => '1',
  6370 => '1',
  6371 => '0',
  6372 => '0',
  6373 => '0',
  6374 => '0',
  6375 => '0',
  6376 => '0',
  6377 => '1',
  6378 => '1',
  6379 => '0',
  6380 => '0',
  6381 => '0',
  6382 => '0',
  6383 => '0',
  6384 => '0',
  6385 => '0',
  6386 => '1',
  6387 => '1',
  6388 => '1',
  6389 => '1',
  6390 => '0',
  6391 => '0',
  6392 => '0',
  6393 => '0',
  6394 => '0',
  6395 => '0',
  6396 => '0',
  6397 => '0',
  6398 => '0',
  6399 => '0',
  6400 => '0',
  6401 => '0',
  6402 => '0',
  6403 => '0',
  6404 => '0',
  6405 => '1',
  6406 => '1',
  6407 => '0',
  6408 => '0',
  6409 => '0',
  6410 => '0',
  6411 => '0',
  6412 => '0',
  6413 => '1',
  6414 => '1',
  6415 => '0',
  6416 => '0',
  6417 => '0',
  6418 => '1',
  6419 => '1',
  6420 => '1',
  6421 => '1',
  6422 => '1',
  6423 => '0',
  6424 => '0',
  6425 => '1',
  6426 => '1',
  6427 => '0',
  6428 => '0',
  6429 => '1',
  6430 => '1',
  6431 => '0',
  6432 => '0',
  6433 => '1',
  6434 => '1',
  6435 => '0',
  6436 => '0',
  6437 => '1',
  6438 => '1',
  6439 => '0',
  6440 => '0',
  6441 => '1',
  6442 => '1',
  6443 => '0',
  6444 => '0',
  6445 => '1',
  6446 => '1',
  6447 => '0',
  6448 => '0',
  6449 => '0',
  6450 => '1',
  6451 => '1',
  6452 => '1',
  6453 => '1',
  6454 => '1',
  6455 => '0',
  6456 => '0',
  6457 => '0',
  6458 => '0',
  6459 => '0',
  6460 => '0',
  6461 => '0',
  6462 => '0',
  6463 => '0',
  6464 => '0',
  6465 => '0',
  6466 => '0',
  6467 => '0',
  6468 => '0',
  6469 => '0',
  6470 => '0',
  6471 => '0',
  6472 => '0',
  6473 => '0',
  6474 => '0',
  6475 => '0',
  6476 => '0',
  6477 => '0',
  6478 => '0',
  6479 => '0',
  6480 => '0',
  6481 => '0',
  6482 => '1',
  6483 => '1',
  6484 => '1',
  6485 => '1',
  6486 => '0',
  6487 => '0',
  6488 => '0',
  6489 => '1',
  6490 => '1',
  6491 => '0',
  6492 => '0',
  6493 => '1',
  6494 => '1',
  6495 => '0',
  6496 => '0',
  6497 => '1',
  6498 => '1',
  6499 => '1',
  6500 => '1',
  6501 => '1',
  6502 => '1',
  6503 => '0',
  6504 => '0',
  6505 => '1',
  6506 => '1',
  6507 => '0',
  6508 => '0',
  6509 => '0',
  6510 => '0',
  6511 => '0',
  6512 => '0',
  6513 => '0',
  6514 => '1',
  6515 => '1',
  6516 => '1',
  6517 => '1',
  6518 => '0',
  6519 => '0',
  6520 => '0',
  6521 => '0',
  6522 => '0',
  6523 => '0',
  6524 => '0',
  6525 => '0',
  6526 => '0',
  6527 => '0',
  6528 => '0',
  6529 => '0',
  6530 => '0',
  6531 => '1',
  6532 => '1',
  6533 => '1',
  6534 => '0',
  6535 => '0',
  6536 => '0',
  6537 => '0',
  6538 => '1',
  6539 => '1',
  6540 => '0',
  6541 => '0',
  6542 => '0',
  6543 => '0',
  6544 => '0',
  6545 => '1',
  6546 => '1',
  6547 => '1',
  6548 => '1',
  6549 => '1',
  6550 => '0',
  6551 => '0',
  6552 => '0',
  6553 => '0',
  6554 => '1',
  6555 => '1',
  6556 => '0',
  6557 => '0',
  6558 => '0',
  6559 => '0',
  6560 => '0',
  6561 => '0',
  6562 => '1',
  6563 => '1',
  6564 => '0',
  6565 => '0',
  6566 => '0',
  6567 => '0',
  6568 => '0',
  6569 => '0',
  6570 => '1',
  6571 => '1',
  6572 => '0',
  6573 => '0',
  6574 => '0',
  6575 => '0',
  6576 => '0',
  6577 => '0',
  6578 => '1',
  6579 => '1',
  6580 => '0',
  6581 => '0',
  6582 => '0',
  6583 => '0',
  6584 => '0',
  6585 => '0',
  6586 => '0',
  6587 => '0',
  6588 => '0',
  6589 => '0',
  6590 => '0',
  6591 => '0',
  6592 => '0',
  6593 => '0',
  6594 => '0',
  6595 => '0',
  6596 => '0',
  6597 => '0',
  6598 => '0',
  6599 => '0',
  6600 => '0',
  6601 => '0',
  6602 => '0',
  6603 => '0',
  6604 => '0',
  6605 => '0',
  6606 => '0',
  6607 => '0',
  6608 => '0',
  6609 => '0',
  6610 => '1',
  6611 => '1',
  6612 => '1',
  6613 => '1',
  6614 => '1',
  6615 => '0',
  6616 => '0',
  6617 => '1',
  6618 => '1',
  6619 => '0',
  6620 => '0',
  6621 => '1',
  6622 => '1',
  6623 => '0',
  6624 => '0',
  6625 => '1',
  6626 => '1',
  6627 => '0',
  6628 => '0',
  6629 => '1',
  6630 => '1',
  6631 => '0',
  6632 => '0',
  6633 => '0',
  6634 => '1',
  6635 => '1',
  6636 => '1',
  6637 => '1',
  6638 => '1',
  6639 => '0',
  6640 => '0',
  6641 => '0',
  6642 => '0',
  6643 => '0',
  6644 => '0',
  6645 => '1',
  6646 => '1',
  6647 => '0',
  6648 => '0',
  6649 => '0',
  6650 => '1',
  6651 => '1',
  6652 => '1',
  6653 => '1',
  6654 => '0',
  6655 => '0',
  6656 => '0',
  6657 => '1',
  6658 => '1',
  6659 => '0',
  6660 => '0',
  6661 => '0',
  6662 => '0',
  6663 => '0',
  6664 => '0',
  6665 => '1',
  6666 => '1',
  6667 => '0',
  6668 => '0',
  6669 => '0',
  6670 => '0',
  6671 => '0',
  6672 => '0',
  6673 => '1',
  6674 => '1',
  6675 => '1',
  6676 => '1',
  6677 => '1',
  6678 => '0',
  6679 => '0',
  6680 => '0',
  6681 => '1',
  6682 => '1',
  6683 => '0',
  6684 => '0',
  6685 => '1',
  6686 => '1',
  6687 => '0',
  6688 => '0',
  6689 => '1',
  6690 => '1',
  6691 => '0',
  6692 => '0',
  6693 => '1',
  6694 => '1',
  6695 => '0',
  6696 => '0',
  6697 => '1',
  6698 => '1',
  6699 => '0',
  6700 => '0',
  6701 => '1',
  6702 => '1',
  6703 => '0',
  6704 => '0',
  6705 => '1',
  6706 => '1',
  6707 => '0',
  6708 => '0',
  6709 => '1',
  6710 => '1',
  6711 => '0',
  6712 => '0',
  6713 => '0',
  6714 => '0',
  6715 => '0',
  6716 => '0',
  6717 => '0',
  6718 => '0',
  6719 => '0',
  6720 => '0',
  6721 => '0',
  6722 => '0',
  6723 => '1',
  6724 => '1',
  6725 => '0',
  6726 => '0',
  6727 => '0',
  6728 => '0',
  6729 => '0',
  6730 => '0',
  6731 => '0',
  6732 => '0',
  6733 => '0',
  6734 => '0',
  6735 => '0',
  6736 => '0',
  6737 => '0',
  6738 => '0',
  6739 => '1',
  6740 => '1',
  6741 => '0',
  6742 => '0',
  6743 => '0',
  6744 => '0',
  6745 => '0',
  6746 => '0',
  6747 => '1',
  6748 => '1',
  6749 => '0',
  6750 => '0',
  6751 => '0',
  6752 => '0',
  6753 => '0',
  6754 => '0',
  6755 => '1',
  6756 => '1',
  6757 => '0',
  6758 => '0',
  6759 => '0',
  6760 => '0',
  6761 => '0',
  6762 => '0',
  6763 => '1',
  6764 => '1',
  6765 => '0',
  6766 => '0',
  6767 => '0',
  6768 => '0',
  6769 => '0',
  6770 => '0',
  6771 => '0',
  6772 => '1',
  6773 => '1',
  6774 => '0',
  6775 => '0',
  6776 => '0',
  6777 => '0',
  6778 => '0',
  6779 => '0',
  6780 => '0',
  6781 => '0',
  6782 => '0',
  6783 => '0',
  6784 => '0',
  6785 => '0',
  6786 => '0',
  6787 => '0',
  6788 => '1',
  6789 => '1',
  6790 => '0',
  6791 => '0',
  6792 => '0',
  6793 => '0',
  6794 => '0',
  6795 => '0',
  6796 => '0',
  6797 => '0',
  6798 => '0',
  6799 => '0',
  6800 => '0',
  6801 => '0',
  6802 => '0',
  6803 => '0',
  6804 => '1',
  6805 => '1',
  6806 => '0',
  6807 => '0',
  6808 => '0',
  6809 => '0',
  6810 => '0',
  6811 => '0',
  6812 => '1',
  6813 => '1',
  6814 => '0',
  6815 => '0',
  6816 => '0',
  6817 => '0',
  6818 => '0',
  6819 => '0',
  6820 => '1',
  6821 => '1',
  6822 => '0',
  6823 => '0',
  6824 => '0',
  6825 => '0',
  6826 => '0',
  6827 => '0',
  6828 => '1',
  6829 => '1',
  6830 => '0',
  6831 => '0',
  6832 => '0',
  6833 => '0',
  6834 => '0',
  6835 => '0',
  6836 => '1',
  6837 => '1',
  6838 => '0',
  6839 => '0',
  6840 => '0',
  6841 => '1',
  6842 => '1',
  6843 => '1',
  6844 => '1',
  6845 => '0',
  6846 => '0',
  6847 => '0',
  6848 => '0',
  6849 => '1',
  6850 => '1',
  6851 => '0',
  6852 => '0',
  6853 => '0',
  6854 => '0',
  6855 => '0',
  6856 => '0',
  6857 => '1',
  6858 => '1',
  6859 => '0',
  6860 => '0',
  6861 => '0',
  6862 => '0',
  6863 => '0',
  6864 => '0',
  6865 => '1',
  6866 => '1',
  6867 => '0',
  6868 => '0',
  6869 => '1',
  6870 => '1',
  6871 => '0',
  6872 => '0',
  6873 => '1',
  6874 => '1',
  6875 => '0',
  6876 => '1',
  6877 => '1',
  6878 => '0',
  6879 => '0',
  6880 => '0',
  6881 => '1',
  6882 => '1',
  6883 => '1',
  6884 => '1',
  6885 => '0',
  6886 => '0',
  6887 => '0',
  6888 => '0',
  6889 => '1',
  6890 => '1',
  6891 => '0',
  6892 => '1',
  6893 => '1',
  6894 => '0',
  6895 => '0',
  6896 => '0',
  6897 => '1',
  6898 => '1',
  6899 => '0',
  6900 => '0',
  6901 => '1',
  6902 => '1',
  6903 => '0',
  6904 => '0',
  6905 => '0',
  6906 => '0',
  6907 => '0',
  6908 => '0',
  6909 => '0',
  6910 => '0',
  6911 => '0',
  6912 => '0',
  6913 => '0',
  6914 => '0',
  6915 => '1',
  6916 => '1',
  6917 => '0',
  6918 => '0',
  6919 => '0',
  6920 => '0',
  6921 => '0',
  6922 => '0',
  6923 => '1',
  6924 => '1',
  6925 => '0',
  6926 => '0',
  6927 => '0',
  6928 => '0',
  6929 => '0',
  6930 => '0',
  6931 => '1',
  6932 => '1',
  6933 => '0',
  6934 => '0',
  6935 => '0',
  6936 => '0',
  6937 => '0',
  6938 => '0',
  6939 => '1',
  6940 => '1',
  6941 => '0',
  6942 => '0',
  6943 => '0',
  6944 => '0',
  6945 => '0',
  6946 => '0',
  6947 => '1',
  6948 => '1',
  6949 => '0',
  6950 => '0',
  6951 => '0',
  6952 => '0',
  6953 => '0',
  6954 => '0',
  6955 => '1',
  6956 => '1',
  6957 => '0',
  6958 => '0',
  6959 => '0',
  6960 => '0',
  6961 => '0',
  6962 => '0',
  6963 => '0',
  6964 => '1',
  6965 => '1',
  6966 => '0',
  6967 => '0',
  6968 => '0',
  6969 => '0',
  6970 => '0',
  6971 => '0',
  6972 => '0',
  6973 => '0',
  6974 => '0',
  6975 => '0',
  6976 => '0',
  6977 => '0',
  6978 => '0',
  6979 => '0',
  6980 => '0',
  6981 => '0',
  6982 => '0',
  6983 => '0',
  6984 => '0',
  6985 => '0',
  6986 => '0',
  6987 => '0',
  6988 => '0',
  6989 => '0',
  6990 => '0',
  6991 => '0',
  6992 => '1',
  6993 => '1',
  6994 => '1',
  6995 => '0',
  6996 => '1',
  6997 => '1',
  6998 => '0',
  6999 => '0',
  7000 => '1',
  7001 => '1',
  7002 => '1',
  7003 => '1',
  7004 => '1',
  7005 => '1',
  7006 => '1',
  7007 => '0',
  7008 => '1',
  7009 => '1',
  7010 => '0',
  7011 => '1',
  7012 => '0',
  7013 => '1',
  7014 => '1',
  7015 => '0',
  7016 => '1',
  7017 => '1',
  7018 => '0',
  7019 => '0',
  7020 => '0',
  7021 => '1',
  7022 => '1',
  7023 => '0',
  7024 => '1',
  7025 => '1',
  7026 => '0',
  7027 => '0',
  7028 => '0',
  7029 => '1',
  7030 => '1',
  7031 => '0',
  7032 => '0',
  7033 => '0',
  7034 => '0',
  7035 => '0',
  7036 => '0',
  7037 => '0',
  7038 => '0',
  7039 => '0',
  7040 => '0',
  7041 => '0',
  7042 => '0',
  7043 => '0',
  7044 => '0',
  7045 => '0',
  7046 => '0',
  7047 => '0',
  7048 => '0',
  7049 => '0',
  7050 => '0',
  7051 => '0',
  7052 => '0',
  7053 => '0',
  7054 => '0',
  7055 => '0',
  7056 => '0',
  7057 => '1',
  7058 => '1',
  7059 => '1',
  7060 => '1',
  7061 => '1',
  7062 => '0',
  7063 => '0',
  7064 => '0',
  7065 => '1',
  7066 => '1',
  7067 => '0',
  7068 => '0',
  7069 => '1',
  7070 => '1',
  7071 => '0',
  7072 => '0',
  7073 => '1',
  7074 => '1',
  7075 => '0',
  7076 => '0',
  7077 => '1',
  7078 => '1',
  7079 => '0',
  7080 => '0',
  7081 => '1',
  7082 => '1',
  7083 => '0',
  7084 => '0',
  7085 => '1',
  7086 => '1',
  7087 => '0',
  7088 => '0',
  7089 => '1',
  7090 => '1',
  7091 => '0',
  7092 => '0',
  7093 => '1',
  7094 => '1',
  7095 => '0',
  7096 => '0',
  7097 => '0',
  7098 => '0',
  7099 => '0',
  7100 => '0',
  7101 => '0',
  7102 => '0',
  7103 => '0',
  7104 => '0',
  7105 => '0',
  7106 => '0',
  7107 => '0',
  7108 => '0',
  7109 => '0',
  7110 => '0',
  7111 => '0',
  7112 => '0',
  7113 => '0',
  7114 => '0',
  7115 => '0',
  7116 => '0',
  7117 => '0',
  7118 => '0',
  7119 => '0',
  7120 => '0',
  7121 => '0',
  7122 => '1',
  7123 => '1',
  7124 => '1',
  7125 => '1',
  7126 => '0',
  7127 => '0',
  7128 => '0',
  7129 => '1',
  7130 => '1',
  7131 => '0',
  7132 => '0',
  7133 => '1',
  7134 => '1',
  7135 => '0',
  7136 => '0',
  7137 => '1',
  7138 => '1',
  7139 => '0',
  7140 => '0',
  7141 => '1',
  7142 => '1',
  7143 => '0',
  7144 => '0',
  7145 => '1',
  7146 => '1',
  7147 => '0',
  7148 => '0',
  7149 => '1',
  7150 => '1',
  7151 => '0',
  7152 => '0',
  7153 => '0',
  7154 => '1',
  7155 => '1',
  7156 => '1',
  7157 => '1',
  7158 => '0',
  7159 => '0',
  7160 => '0',
  7161 => '0',
  7162 => '0',
  7163 => '0',
  7164 => '0',
  7165 => '0',
  7166 => '0',
  7167 => '0',
  7168 => '0',
  7169 => '0',
  7170 => '0',
  7171 => '0',
  7172 => '0',
  7173 => '0',
  7174 => '0',
  7175 => '0',
  7176 => '0',
  7177 => '0',
  7178 => '0',
  7179 => '0',
  7180 => '0',
  7181 => '0',
  7182 => '0',
  7183 => '0',
  7184 => '0',
  7185 => '1',
  7186 => '1',
  7187 => '1',
  7188 => '1',
  7189 => '1',
  7190 => '0',
  7191 => '0',
  7192 => '0',
  7193 => '1',
  7194 => '1',
  7195 => '0',
  7196 => '0',
  7197 => '1',
  7198 => '1',
  7199 => '0',
  7200 => '0',
  7201 => '1',
  7202 => '1',
  7203 => '0',
  7204 => '0',
  7205 => '1',
  7206 => '1',
  7207 => '0',
  7208 => '0',
  7209 => '1',
  7210 => '1',
  7211 => '1',
  7212 => '1',
  7213 => '1',
  7214 => '0',
  7215 => '0',
  7216 => '0',
  7217 => '1',
  7218 => '1',
  7219 => '0',
  7220 => '0',
  7221 => '0',
  7222 => '0',
  7223 => '0',
  7224 => '0',
  7225 => '1',
  7226 => '1',
  7227 => '0',
  7228 => '0',
  7229 => '0',
  7230 => '0',
  7231 => '0',
  7232 => '0',
  7233 => '0',
  7234 => '0',
  7235 => '0',
  7236 => '0',
  7237 => '0',
  7238 => '0',
  7239 => '0',
  7240 => '0',
  7241 => '0',
  7242 => '0',
  7243 => '0',
  7244 => '0',
  7245 => '0',
  7246 => '0',
  7247 => '0',
  7248 => '0',
  7249 => '0',
  7250 => '1',
  7251 => '1',
  7252 => '1',
  7253 => '1',
  7254 => '1',
  7255 => '0',
  7256 => '0',
  7257 => '1',
  7258 => '1',
  7259 => '0',
  7260 => '0',
  7261 => '1',
  7262 => '1',
  7263 => '0',
  7264 => '0',
  7265 => '1',
  7266 => '1',
  7267 => '0',
  7268 => '0',
  7269 => '1',
  7270 => '1',
  7271 => '0',
  7272 => '0',
  7273 => '0',
  7274 => '1',
  7275 => '1',
  7276 => '1',
  7277 => '1',
  7278 => '1',
  7279 => '0',
  7280 => '0',
  7281 => '0',
  7282 => '0',
  7283 => '0',
  7284 => '0',
  7285 => '1',
  7286 => '1',
  7287 => '0',
  7288 => '0',
  7289 => '0',
  7290 => '0',
  7291 => '0',
  7292 => '0',
  7293 => '1',
  7294 => '1',
  7295 => '0',
  7296 => '0',
  7297 => '0',
  7298 => '0',
  7299 => '0',
  7300 => '0',
  7301 => '0',
  7302 => '0',
  7303 => '0',
  7304 => '0',
  7305 => '0',
  7306 => '0',
  7307 => '0',
  7308 => '0',
  7309 => '0',
  7310 => '0',
  7311 => '0',
  7312 => '0',
  7313 => '1',
  7314 => '1',
  7315 => '1',
  7316 => '1',
  7317 => '1',
  7318 => '0',
  7319 => '0',
  7320 => '0',
  7321 => '1',
  7322 => '1',
  7323 => '0',
  7324 => '0',
  7325 => '1',
  7326 => '1',
  7327 => '0',
  7328 => '0',
  7329 => '1',
  7330 => '1',
  7331 => '0',
  7332 => '0',
  7333 => '0',
  7334 => '0',
  7335 => '0',
  7336 => '0',
  7337 => '1',
  7338 => '1',
  7339 => '0',
  7340 => '0',
  7341 => '0',
  7342 => '0',
  7343 => '0',
  7344 => '0',
  7345 => '1',
  7346 => '1',
  7347 => '0',
  7348 => '0',
  7349 => '0',
  7350 => '0',
  7351 => '0',
  7352 => '0',
  7353 => '0',
  7354 => '0',
  7355 => '0',
  7356 => '0',
  7357 => '0',
  7358 => '0',
  7359 => '0',
  7360 => '0',
  7361 => '0',
  7362 => '0',
  7363 => '0',
  7364 => '0',
  7365 => '0',
  7366 => '0',
  7367 => '0',
  7368 => '0',
  7369 => '0',
  7370 => '0',
  7371 => '0',
  7372 => '0',
  7373 => '0',
  7374 => '0',
  7375 => '0',
  7376 => '0',
  7377 => '0',
  7378 => '1',
  7379 => '1',
  7380 => '1',
  7381 => '1',
  7382 => '0',
  7383 => '0',
  7384 => '0',
  7385 => '1',
  7386 => '1',
  7387 => '0',
  7388 => '0',
  7389 => '0',
  7390 => '0',
  7391 => '0',
  7392 => '0',
  7393 => '0',
  7394 => '1',
  7395 => '1',
  7396 => '1',
  7397 => '1',
  7398 => '0',
  7399 => '0',
  7400 => '0',
  7401 => '0',
  7402 => '0',
  7403 => '0',
  7404 => '0',
  7405 => '1',
  7406 => '1',
  7407 => '0',
  7408 => '0',
  7409 => '1',
  7410 => '1',
  7411 => '1',
  7412 => '1',
  7413 => '1',
  7414 => '0',
  7415 => '0',
  7416 => '0',
  7417 => '0',
  7418 => '0',
  7419 => '0',
  7420 => '0',
  7421 => '0',
  7422 => '0',
  7423 => '0',
  7424 => '0',
  7425 => '0',
  7426 => '1',
  7427 => '1',
  7428 => '0',
  7429 => '0',
  7430 => '0',
  7431 => '0',
  7432 => '0',
  7433 => '0',
  7434 => '1',
  7435 => '1',
  7436 => '0',
  7437 => '0',
  7438 => '0',
  7439 => '0',
  7440 => '0',
  7441 => '1',
  7442 => '1',
  7443 => '1',
  7444 => '1',
  7445 => '1',
  7446 => '0',
  7447 => '0',
  7448 => '0',
  7449 => '0',
  7450 => '1',
  7451 => '1',
  7452 => '0',
  7453 => '0',
  7454 => '0',
  7455 => '0',
  7456 => '0',
  7457 => '0',
  7458 => '1',
  7459 => '1',
  7460 => '0',
  7461 => '0',
  7462 => '0',
  7463 => '0',
  7464 => '0',
  7465 => '0',
  7466 => '1',
  7467 => '1',
  7468 => '0',
  7469 => '0',
  7470 => '0',
  7471 => '0',
  7472 => '0',
  7473 => '0',
  7474 => '0',
  7475 => '1',
  7476 => '1',
  7477 => '1',
  7478 => '0',
  7479 => '0',
  7480 => '0',
  7481 => '0',
  7482 => '0',
  7483 => '0',
  7484 => '0',
  7485 => '0',
  7486 => '0',
  7487 => '0',
  7488 => '0',
  7489 => '0',
  7490 => '0',
  7491 => '0',
  7492 => '0',
  7493 => '0',
  7494 => '0',
  7495 => '0',
  7496 => '0',
  7497 => '0',
  7498 => '0',
  7499 => '0',
  7500 => '0',
  7501 => '0',
  7502 => '0',
  7503 => '0',
  7504 => '0',
  7505 => '1',
  7506 => '1',
  7507 => '0',
  7508 => '0',
  7509 => '1',
  7510 => '1',
  7511 => '0',
  7512 => '0',
  7513 => '1',
  7514 => '1',
  7515 => '0',
  7516 => '0',
  7517 => '1',
  7518 => '1',
  7519 => '0',
  7520 => '0',
  7521 => '1',
  7522 => '1',
  7523 => '0',
  7524 => '0',
  7525 => '1',
  7526 => '1',
  7527 => '0',
  7528 => '0',
  7529 => '1',
  7530 => '1',
  7531 => '0',
  7532 => '0',
  7533 => '1',
  7534 => '1',
  7535 => '0',
  7536 => '0',
  7537 => '0',
  7538 => '1',
  7539 => '1',
  7540 => '1',
  7541 => '1',
  7542 => '1',
  7543 => '0',
  7544 => '0',
  7545 => '0',
  7546 => '0',
  7547 => '0',
  7548 => '0',
  7549 => '0',
  7550 => '0',
  7551 => '0',
  7552 => '0',
  7553 => '0',
  7554 => '0',
  7555 => '0',
  7556 => '0',
  7557 => '0',
  7558 => '0',
  7559 => '0',
  7560 => '0',
  7561 => '0',
  7562 => '0',
  7563 => '0',
  7564 => '0',
  7565 => '0',
  7566 => '0',
  7567 => '0',
  7568 => '0',
  7569 => '1',
  7570 => '1',
  7571 => '0',
  7572 => '0',
  7573 => '1',
  7574 => '1',
  7575 => '0',
  7576 => '0',
  7577 => '1',
  7578 => '1',
  7579 => '0',
  7580 => '0',
  7581 => '1',
  7582 => '1',
  7583 => '0',
  7584 => '0',
  7585 => '1',
  7586 => '1',
  7587 => '0',
  7588 => '0',
  7589 => '1',
  7590 => '1',
  7591 => '0',
  7592 => '0',
  7593 => '0',
  7594 => '1',
  7595 => '1',
  7596 => '1',
  7597 => '1',
  7598 => '0',
  7599 => '0',
  7600 => '0',
  7601 => '0',
  7602 => '0',
  7603 => '1',
  7604 => '1',
  7605 => '0',
  7606 => '0',
  7607 => '0',
  7608 => '0',
  7609 => '0',
  7610 => '0',
  7611 => '0',
  7612 => '0',
  7613 => '0',
  7614 => '0',
  7615 => '0',
  7616 => '0',
  7617 => '0',
  7618 => '0',
  7619 => '0',
  7620 => '0',
  7621 => '0',
  7622 => '0',
  7623 => '0',
  7624 => '0',
  7625 => '0',
  7626 => '0',
  7627 => '0',
  7628 => '0',
  7629 => '0',
  7630 => '0',
  7631 => '0',
  7632 => '1',
  7633 => '1',
  7634 => '0',
  7635 => '0',
  7636 => '0',
  7637 => '1',
  7638 => '1',
  7639 => '0',
  7640 => '1',
  7641 => '1',
  7642 => '0',
  7643 => '0',
  7644 => '0',
  7645 => '1',
  7646 => '1',
  7647 => '0',
  7648 => '1',
  7649 => '1',
  7650 => '0',
  7651 => '1',
  7652 => '0',
  7653 => '1',
  7654 => '1',
  7655 => '0',
  7656 => '1',
  7657 => '1',
  7658 => '1',
  7659 => '1',
  7660 => '1',
  7661 => '1',
  7662 => '1',
  7663 => '0',
  7664 => '0',
  7665 => '1',
  7666 => '1',
  7667 => '0',
  7668 => '1',
  7669 => '1',
  7670 => '0',
  7671 => '0',
  7672 => '0',
  7673 => '0',
  7674 => '0',
  7675 => '0',
  7676 => '0',
  7677 => '0',
  7678 => '0',
  7679 => '0',
  7680 => '0',
  7681 => '0',
  7682 => '0',
  7683 => '0',
  7684 => '0',
  7685 => '0',
  7686 => '0',
  7687 => '0',
  7688 => '0',
  7689 => '0',
  7690 => '0',
  7691 => '0',
  7692 => '0',
  7693 => '0',
  7694 => '0',
  7695 => '0',
  7696 => '1',
  7697 => '1',
  7698 => '0',
  7699 => '0',
  7700 => '0',
  7701 => '1',
  7702 => '1',
  7703 => '0',
  7704 => '0',
  7705 => '1',
  7706 => '1',
  7707 => '0',
  7708 => '1',
  7709 => '1',
  7710 => '0',
  7711 => '0',
  7712 => '0',
  7713 => '0',
  7714 => '1',
  7715 => '1',
  7716 => '1',
  7717 => '0',
  7718 => '0',
  7719 => '0',
  7720 => '0',
  7721 => '1',
  7722 => '1',
  7723 => '0',
  7724 => '1',
  7725 => '1',
  7726 => '0',
  7727 => '0',
  7728 => '1',
  7729 => '1',
  7730 => '0',
  7731 => '0',
  7732 => '0',
  7733 => '1',
  7734 => '1',
  7735 => '0',
  7736 => '0',
  7737 => '0',
  7738 => '0',
  7739 => '0',
  7740 => '0',
  7741 => '0',
  7742 => '0',
  7743 => '0',
  7744 => '0',
  7745 => '0',
  7746 => '0',
  7747 => '0',
  7748 => '0',
  7749 => '0',
  7750 => '0',
  7751 => '0',
  7752 => '0',
  7753 => '0',
  7754 => '0',
  7755 => '0',
  7756 => '0',
  7757 => '0',
  7758 => '0',
  7759 => '0',
  7760 => '0',
  7761 => '1',
  7762 => '1',
  7763 => '0',
  7764 => '0',
  7765 => '1',
  7766 => '1',
  7767 => '0',
  7768 => '0',
  7769 => '1',
  7770 => '1',
  7771 => '0',
  7772 => '0',
  7773 => '1',
  7774 => '1',
  7775 => '0',
  7776 => '0',
  7777 => '1',
  7778 => '1',
  7779 => '0',
  7780 => '0',
  7781 => '1',
  7782 => '1',
  7783 => '0',
  7784 => '0',
  7785 => '0',
  7786 => '1',
  7787 => '1',
  7788 => '1',
  7789 => '1',
  7790 => '0',
  7791 => '0',
  7792 => '0',
  7793 => '0',
  7794 => '0',
  7795 => '1',
  7796 => '1',
  7797 => '0',
  7798 => '0',
  7799 => '0',
  7800 => '0',
  7801 => '0',
  7802 => '1',
  7803 => '1',
  7804 => '0',
  7805 => '0',
  7806 => '0',
  7807 => '0',
  7808 => '0',
  7809 => '0',
  7810 => '0',
  7811 => '0',
  7812 => '0',
  7813 => '0',
  7814 => '0',
  7815 => '0',
  7816 => '0',
  7817 => '0',
  7818 => '0',
  7819 => '0',
  7820 => '0',
  7821 => '0',
  7822 => '0',
  7823 => '0',
  7824 => '0',
  7825 => '1',
  7826 => '1',
  7827 => '1',
  7828 => '1',
  7829 => '1',
  7830 => '1',
  7831 => '0',
  7832 => '0',
  7833 => '0',
  7834 => '0',
  7835 => '0',
  7836 => '1',
  7837 => '1',
  7838 => '0',
  7839 => '0',
  7840 => '0',
  7841 => '0',
  7842 => '0',
  7843 => '1',
  7844 => '1',
  7845 => '0',
  7846 => '0',
  7847 => '0',
  7848 => '0',
  7849 => '0',
  7850 => '1',
  7851 => '1',
  7852 => '0',
  7853 => '0',
  7854 => '0',
  7855 => '0',
  7856 => '0',
  7857 => '1',
  7858 => '1',
  7859 => '1',
  7860 => '1',
  7861 => '1',
  7862 => '1',
  7863 => '0',
  7864 => '0',
  7865 => '0',
  7866 => '0',
  7867 => '0',
  7868 => '0',
  7869 => '0',
  7870 => '0',
  7871 => '0',
  7872 => '0',
  7873 => '0',
  7874 => '0',
  7875 => '0',
  7876 => '1',
  7877 => '1',
  7878 => '1',
  7879 => '0',
  7880 => '0',
  7881 => '0',
  7882 => '0',
  7883 => '1',
  7884 => '1',
  7885 => '0',
  7886 => '0',
  7887 => '0',
  7888 => '0',
  7889 => '0',
  7890 => '0',
  7891 => '1',
  7892 => '1',
  7893 => '0',
  7894 => '0',
  7895 => '0',
  7896 => '0',
  7897 => '1',
  7898 => '1',
  7899 => '1',
  7900 => '0',
  7901 => '0',
  7902 => '0',
  7903 => '0',
  7904 => '0',
  7905 => '0',
  7906 => '0',
  7907 => '1',
  7908 => '1',
  7909 => '0',
  7910 => '0',
  7911 => '0',
  7912 => '0',
  7913 => '0',
  7914 => '0',
  7915 => '1',
  7916 => '1',
  7917 => '0',
  7918 => '0',
  7919 => '0',
  7920 => '0',
  7921 => '0',
  7922 => '0',
  7923 => '0',
  7924 => '1',
  7925 => '1',
  7926 => '1',
  7927 => '0',
  7928 => '0',
  7929 => '0',
  7930 => '0',
  7931 => '0',
  7932 => '0',
  7933 => '0',
  7934 => '0',
  7935 => '0',
  7936 => '0',
  7937 => '0',
  7938 => '0',
  7939 => '1',
  7940 => '1',
  7941 => '0',
  7942 => '0',
  7943 => '0',
  7944 => '0',
  7945 => '0',
  7946 => '0',
  7947 => '1',
  7948 => '1',
  7949 => '0',
  7950 => '0',
  7951 => '0',
  7952 => '0',
  7953 => '0',
  7954 => '0',
  7955 => '1',
  7956 => '1',
  7957 => '0',
  7958 => '0',
  7959 => '0',
  7960 => '0',
  7961 => '0',
  7962 => '0',
  7963 => '1',
  7964 => '1',
  7965 => '0',
  7966 => '0',
  7967 => '0',
  7968 => '0',
  7969 => '0',
  7970 => '0',
  7971 => '1',
  7972 => '1',
  7973 => '0',
  7974 => '0',
  7975 => '0',
  7976 => '0',
  7977 => '0',
  7978 => '0',
  7979 => '1',
  7980 => '1',
  7981 => '0',
  7982 => '0',
  7983 => '0',
  7984 => '0',
  7985 => '0',
  7986 => '0',
  7987 => '1',
  7988 => '1',
  7989 => '0',
  7990 => '0',
  7991 => '0',
  7992 => '0',
  7993 => '0',
  7994 => '0',
  7995 => '0',
  7996 => '0',
  7997 => '0',
  7998 => '0',
  7999 => '0',
  8000 => '0',
  8001 => '1',
  8002 => '1',
  8003 => '1',
  8004 => '0',
  8005 => '0',
  8006 => '0',
  8007 => '0',
  8008 => '0',
  8009 => '0',
  8010 => '0',
  8011 => '1',
  8012 => '1',
  8013 => '0',
  8014 => '0',
  8015 => '0',
  8016 => '0',
  8017 => '0',
  8018 => '0',
  8019 => '1',
  8020 => '1',
  8021 => '0',
  8022 => '0',
  8023 => '0',
  8024 => '0',
  8025 => '0',
  8026 => '0',
  8027 => '0',
  8028 => '1',
  8029 => '1',
  8030 => '1',
  8031 => '0',
  8032 => '0',
  8033 => '0',
  8034 => '0',
  8035 => '1',
  8036 => '1',
  8037 => '0',
  8038 => '0',
  8039 => '0',
  8040 => '0',
  8041 => '0',
  8042 => '0',
  8043 => '1',
  8044 => '1',
  8045 => '0',
  8046 => '0',
  8047 => '0',
  8048 => '0',
  8049 => '1',
  8050 => '1',
  8051 => '1',
  8052 => '0',
  8053 => '0',
  8054 => '0',
  8055 => '0',
  8056 => '0',
  8057 => '0',
  8058 => '0',
  8059 => '0',
  8060 => '0',
  8061 => '0',
  8062 => '0',
  8063 => '0',
  8064 => '0',
  8065 => '1',
  8066 => '1',
  8067 => '1',
  8068 => '0',
  8069 => '0',
  8070 => '1',
  8071 => '0',
  8072 => '1',
  8073 => '0',
  8074 => '0',
  8075 => '1',
  8076 => '1',
  8077 => '1',
  8078 => '0',
  8079 => '0',
  8080 => '0',
  8081 => '0',
  8082 => '0',
  8083 => '0',
  8084 => '0',
  8085 => '0',
  8086 => '0',
  8087 => '0',
  8088 => '0',
  8089 => '0',
  8090 => '0',
  8091 => '0',
  8092 => '0',
  8093 => '0',
  8094 => '0',
  8095 => '0',
  8096 => '0',
  8097 => '0',
  8098 => '0',
  8099 => '0',
  8100 => '0',
  8101 => '0',
  8102 => '0',
  8103 => '0',
  8104 => '0',
  8105 => '0',
  8106 => '0',
  8107 => '0',
  8108 => '0',
  8109 => '0',
  8110 => '0',
  8111 => '0',
  8112 => '0',
  8113 => '0',
  8114 => '0',
  8115 => '0',
  8116 => '0',
  8117 => '0',
  8118 => '0',
  8119 => '0',
  8120 => '0',
  8121 => '0',
  8122 => '0',
  8123 => '0',
  8124 => '0',
  8125 => '0',
  8126 => '0',
  8127 => '0',
  8128 => '1',
  8129 => '1',
  8130 => '1',
  8131 => '1',
  8132 => '1',
  8133 => '1',
  8134 => '1',
  8135 => '0',
  8136 => '1',
  8137 => '1',
  8138 => '1',
  8139 => '1',
  8140 => '1',
  8141 => '1',
  8142 => '1',
  8143 => '0',
  8144 => '1',
  8145 => '1',
  8146 => '1',
  8147 => '1',
  8148 => '1',
  8149 => '1',
  8150 => '1',
  8151 => '0',
  8152 => '1',
  8153 => '1',
  8154 => '1',
  8155 => '1',
  8156 => '1',
  8157 => '1',
  8158 => '1',
  8159 => '0',
  8160 => '1',
  8161 => '1',
  8162 => '1',
  8163 => '1',
  8164 => '1',
  8165 => '1',
  8166 => '1',
  8167 => '0',
  8168 => '1',
  8169 => '1',
  8170 => '1',
  8171 => '1',
  8172 => '1',
  8173 => '1',
  8174 => '1',
  8175 => '0',
  8176 => '1',
  8177 => '1',
  8178 => '1',
  8179 => '1',
  8180 => '1',
  8181 => '1',
  8182 => '1',
  8183 => '0',
  8184 => '0',
  8185 => '0',
  8186 => '0',
  8187 => '0',
  8188 => '0',
  8189 => '0',
  8190 => '0',
  8191 => '0',
	others => '0'
);

begin

process (clock)
begin
	if (clock'event and clock = '1') then
		q <= rom(to_integer(unsigned(address(addrbits-1 downto 0))));
	end if;
end process;

end arch;

