-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b0bb5",
     9 => x"a0080b0b",
    10 => x"0bb5a408",
    11 => x"0b0b0bb5",
    12 => x"a8080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"b5a80c0b",
    16 => x"0b0bb5a4",
    17 => x"0c0b0b0b",
    18 => x"b5a00c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0babe4",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"b5a070bb",
    57 => x"d0278b38",
    58 => x"80717084",
    59 => x"05530c81",
    60 => x"e2048c51",
    61 => x"8af10402",
    62 => x"fc050df8",
    63 => x"80518f0b",
    64 => x"b5b00c9f",
    65 => x"0bb5b40c",
    66 => x"a0717081",
    67 => x"055334b5",
    68 => x"b408ff05",
    69 => x"b5b40cb5",
    70 => x"b4088025",
    71 => x"eb38b5b0",
    72 => x"08ff05b5",
    73 => x"b00cb5b0",
    74 => x"088025d7",
    75 => x"38028405",
    76 => x"0d0402f0",
    77 => x"050df880",
    78 => x"53f8a054",
    79 => x"83bf5273",
    80 => x"70810555",
    81 => x"33517073",
    82 => x"70810555",
    83 => x"34ff1252",
    84 => x"718025eb",
    85 => x"38fbc053",
    86 => x"9f52a073",
    87 => x"70810555",
    88 => x"34ff1252",
    89 => x"718025f2",
    90 => x"38029005",
    91 => x"0d0402f4",
    92 => x"050d7453",
    93 => x"8e0bb5b0",
    94 => x"08258f38",
    95 => x"82b22db5",
    96 => x"b008ff05",
    97 => x"b5b00c82",
    98 => x"f404b5b0",
    99 => x"08b5b408",
   100 => x"5351728a",
   101 => x"2e098106",
   102 => x"b7387151",
   103 => x"719f24a0",
   104 => x"38b5b008",
   105 => x"a02911f8",
   106 => x"80115151",
   107 => x"a07134b5",
   108 => x"b4088105",
   109 => x"b5b40cb5",
   110 => x"b408519f",
   111 => x"7125e238",
   112 => x"800bb5b4",
   113 => x"0cb5b008",
   114 => x"8105b5b0",
   115 => x"0c83e404",
   116 => x"70a02912",
   117 => x"f8801151",
   118 => x"51727134",
   119 => x"b5b40881",
   120 => x"05b5b40c",
   121 => x"b5b408a0",
   122 => x"2e098106",
   123 => x"8e38800b",
   124 => x"b5b40cb5",
   125 => x"b0088105",
   126 => x"b5b00c02",
   127 => x"8c050d04",
   128 => x"02e8050d",
   129 => x"77795656",
   130 => x"880bfc16",
   131 => x"77712c8f",
   132 => x"06545254",
   133 => x"80537272",
   134 => x"25953871",
   135 => x"53fbe014",
   136 => x"51877134",
   137 => x"8114ff14",
   138 => x"545472f1",
   139 => x"387153f9",
   140 => x"1576712c",
   141 => x"87065351",
   142 => x"71802e8b",
   143 => x"38fbe014",
   144 => x"51717134",
   145 => x"81145472",
   146 => x"8e249538",
   147 => x"8f733153",
   148 => x"fbe01451",
   149 => x"a0713481",
   150 => x"14ff1454",
   151 => x"5472f138",
   152 => x"0298050d",
   153 => x"0402ec05",
   154 => x"0d800bb5",
   155 => x"b80cf68c",
   156 => x"08f69008",
   157 => x"71882c56",
   158 => x"5481ff06",
   159 => x"52737225",
   160 => x"88387154",
   161 => x"820bb5b8",
   162 => x"0c72882c",
   163 => x"7381ff06",
   164 => x"54557473",
   165 => x"258b3872",
   166 => x"b5b80884",
   167 => x"07b5b80c",
   168 => x"5573842b",
   169 => x"86a07125",
   170 => x"83713170",
   171 => x"0b0b0bb2",
   172 => x"f80c8171",
   173 => x"2bff05f6",
   174 => x"880cfecc",
   175 => x"13ff122c",
   176 => x"788829ff",
   177 => x"94057081",
   178 => x"2cb5b808",
   179 => x"52585255",
   180 => x"51525476",
   181 => x"802e8538",
   182 => x"70810751",
   183 => x"70f6940c",
   184 => x"71098105",
   185 => x"f6800c72",
   186 => x"098105f6",
   187 => x"840c0294",
   188 => x"050d0402",
   189 => x"f4050d74",
   190 => x"53727081",
   191 => x"055480f5",
   192 => x"2d527180",
   193 => x"2e893871",
   194 => x"5182ee2d",
   195 => x"85f90402",
   196 => x"8c050d04",
   197 => x"02f8050d",
   198 => x"a5bd2d80",
   199 => x"da51a6f4",
   200 => x"2db5a008",
   201 => x"812a7081",
   202 => x"06515271",
   203 => x"802ee938",
   204 => x"0288050d",
   205 => x"0402f405",
   206 => x"0dbbc008",
   207 => x"81c406b4",
   208 => x"940b80f5",
   209 => x"2d525270",
   210 => x"802e8638",
   211 => x"71848007",
   212 => x"52b3cc0b",
   213 => x"80f52d72",
   214 => x"07b3e40b",
   215 => x"80f52d70",
   216 => x"812a7081",
   217 => x"06515354",
   218 => x"5270802e",
   219 => x"86387182",
   220 => x"80075272",
   221 => x"81065170",
   222 => x"802e8538",
   223 => x"71880752",
   224 => x"b3f00b80",
   225 => x"f52d7084",
   226 => x"2b730781",
   227 => x"8432b5a0",
   228 => x"0c51028c",
   229 => x"050d0402",
   230 => x"f4050d74",
   231 => x"70818432",
   232 => x"bbc00c70",
   233 => x"83065253",
   234 => x"70b3c40b",
   235 => x"880581b7",
   236 => x"2d72892a",
   237 => x"70810651",
   238 => x"5170b494",
   239 => x"0b81b72d",
   240 => x"72832a81",
   241 => x"0673882a",
   242 => x"70810651",
   243 => x"52527080",
   244 => x"2e853871",
   245 => x"82075271",
   246 => x"b3e40b81",
   247 => x"b72d7284",
   248 => x"2c708306",
   249 => x"515170b3",
   250 => x"f00b81b7",
   251 => x"2d70b5a0",
   252 => x"0c028c05",
   253 => x"0d0402d4",
   254 => x"050daebc",
   255 => x"5185f32d",
   256 => x"9bfb2db5",
   257 => x"a008802e",
   258 => x"82ab3886",
   259 => x"b52db5a0",
   260 => x"08538ed6",
   261 => x"2db5a008",
   262 => x"54b5a008",
   263 => x"802e8297",
   264 => x"389ebe2d",
   265 => x"b5a00880",
   266 => x"2e8738ae",
   267 => x"d45188be",
   268 => x"0497dd2d",
   269 => x"b5a00880",
   270 => x"2e9c38af",
   271 => x"945185f3",
   272 => x"2d86942d",
   273 => x"72840753",
   274 => x"810bfec4",
   275 => x"0c72fec0",
   276 => x"0c725187",
   277 => x"972d840b",
   278 => x"fec40caf",
   279 => x"dc5185f3",
   280 => x"2daff452",
   281 => x"b5c05194",
   282 => x"f22db5a0",
   283 => x"089838b0",
   284 => x"805185f3",
   285 => x"2db09852",
   286 => x"b5c05194",
   287 => x"f22db5a0",
   288 => x"08802e81",
   289 => x"b038b0a4",
   290 => x"5185f32d",
   291 => x"b5c40857",
   292 => x"8077595a",
   293 => x"767a2e8b",
   294 => x"38811a78",
   295 => x"812a595a",
   296 => x"77f738f7",
   297 => x"1a5a8077",
   298 => x"25818038",
   299 => x"79527751",
   300 => x"84802db5",
   301 => x"cc52b5c0",
   302 => x"5197b72d",
   303 => x"b5a00853",
   304 => x"b5a00880",
   305 => x"2e80c938",
   306 => x"b5cc5b80",
   307 => x"5989fd04",
   308 => x"7a708405",
   309 => x"5c087081",
   310 => x"ff067188",
   311 => x"2c7081ff",
   312 => x"0673902c",
   313 => x"7081ff06",
   314 => x"75982afe",
   315 => x"c80cfec8",
   316 => x"0c58fec8",
   317 => x"0c57fec8",
   318 => x"0c841a5a",
   319 => x"53765384",
   320 => x"80772584",
   321 => x"38848053",
   322 => x"727924c4",
   323 => x"388a9b04",
   324 => x"b0c05185",
   325 => x"f32d7254",
   326 => x"8ab704b5",
   327 => x"c051978a",
   328 => x"2dfc8017",
   329 => x"81195957",
   330 => x"89a60482",
   331 => x"0bfec40c",
   332 => x"81548ab7",
   333 => x"04805473",
   334 => x"b5a00c02",
   335 => x"ac050d04",
   336 => x"02f8050d",
   337 => x"a7c42d81",
   338 => x"f72d8151",
   339 => x"84e52dfe",
   340 => x"c4528172",
   341 => x"0ca5852d",
   342 => x"a5852d84",
   343 => x"720c87f6",
   344 => x"2db2fc51",
   345 => x"a8dd2d80",
   346 => x"5184e52d",
   347 => x"0288050d",
   348 => x"0402cc05",
   349 => x"0d8cb851",
   350 => x"87972d81",
   351 => x"0bfec40c",
   352 => x"8cb80bfe",
   353 => x"c00c840b",
   354 => x"fec40ca5",
   355 => x"a02da7b8",
   356 => x"2da5852d",
   357 => x"a5852d81",
   358 => x"f72d8151",
   359 => x"84e52da5",
   360 => x"852da585",
   361 => x"2d815184",
   362 => x"e52dbae8",
   363 => x"51a2cd2d",
   364 => x"b5a008ff",
   365 => x"24f43881",
   366 => x"f452bb90",
   367 => x"51a3912d",
   368 => x"87f62db5",
   369 => x"a008802e",
   370 => x"82b93880",
   371 => x"70715b58",
   372 => x"56947652",
   373 => x"5884e52d",
   374 => x"b2fc51a8",
   375 => x"dd2da585",
   376 => x"2d02b405",
   377 => x"79842905",
   378 => x"f011bae8",
   379 => x"535153a2",
   380 => x"cd2db5a0",
   381 => x"08730cb5",
   382 => x"a008ff2e",
   383 => x"0981068d",
   384 => x"38ff1858",
   385 => x"7780d438",
   386 => x"77598cdb",
   387 => x"04811959",
   388 => x"94587883",
   389 => x"2e098106",
   390 => x"80c13880",
   391 => x"7a8306fe",
   392 => x"cc0c7a70",
   393 => x"852a7081",
   394 => x"067f5851",
   395 => x"55565972",
   396 => x"792e8a38",
   397 => x"73fe8032",
   398 => x"16568cc0",
   399 => x"04731656",
   400 => x"74842a70",
   401 => x"81067c56",
   402 => x"51537280",
   403 => x"2e8a3873",
   404 => x"fe803217",
   405 => x"578cdb04",
   406 => x"73175776",
   407 => x"76075372",
   408 => x"802e80d0",
   409 => x"38fed008",
   410 => x"70810651",
   411 => x"5372802e",
   412 => x"80c23876",
   413 => x"76555380",
   414 => x"ff772584",
   415 => x"3880ff53",
   416 => x"80ff7425",
   417 => x"843880ff",
   418 => x"5472ff80",
   419 => x"258438ff",
   420 => x"805373ff",
   421 => x"80258438",
   422 => x"ff805476",
   423 => x"73317675",
   424 => x"3174882b",
   425 => x"83fe8006",
   426 => x"7681ff06",
   427 => x"7107fed0",
   428 => x"0c555757",
   429 => x"a5bd2da8",
   430 => x"ed2db5a0",
   431 => x"085486b5",
   432 => x"2db5a008",
   433 => x"fec00c86",
   434 => x"b52db5a0",
   435 => x"08b5bc08",
   436 => x"2e9c38b5",
   437 => x"a008b5bc",
   438 => x"0c845373",
   439 => x"5184e52d",
   440 => x"a5852da5",
   441 => x"852dff13",
   442 => x"53728025",
   443 => x"ee387380",
   444 => x"2e89388a",
   445 => x"0bfec40c",
   446 => x"8bde0482",
   447 => x"0bfec40c",
   448 => x"8bde04b0",
   449 => x"d45185f3",
   450 => x"2d820bfe",
   451 => x"c40c800b",
   452 => x"b5a00c02",
   453 => x"b4050d04",
   454 => x"02e8050d",
   455 => x"77797b58",
   456 => x"55558053",
   457 => x"727625a3",
   458 => x"38747081",
   459 => x"055680f5",
   460 => x"2d747081",
   461 => x"055680f5",
   462 => x"2d525271",
   463 => x"712e8638",
   464 => x"81518ecd",
   465 => x"04811353",
   466 => x"8ea40480",
   467 => x"5170b5a0",
   468 => x"0c029805",
   469 => x"0d0402d8",
   470 => x"050d800b",
   471 => x"b9d40cb5",
   472 => x"cc528051",
   473 => x"9d9b2db5",
   474 => x"a00854b5",
   475 => x"a0088c38",
   476 => x"b0ec5185",
   477 => x"f32d7355",
   478 => x"93fb0480",
   479 => x"56810bb9",
   480 => x"f80c8853",
   481 => x"b18052b6",
   482 => x"82518e98",
   483 => x"2db5a008",
   484 => x"762e0981",
   485 => x"068738b5",
   486 => x"a008b9f8",
   487 => x"0c8853b1",
   488 => x"8c52b69e",
   489 => x"518e982d",
   490 => x"b5a00887",
   491 => x"38b5a008",
   492 => x"b9f80cb9",
   493 => x"f80852b1",
   494 => x"9851a0b8",
   495 => x"2db9f808",
   496 => x"802e80f6",
   497 => x"38b9920b",
   498 => x"80f52db9",
   499 => x"930b80f5",
   500 => x"2d71982b",
   501 => x"71902b07",
   502 => x"b9940b80",
   503 => x"f52d7088",
   504 => x"2b7207b9",
   505 => x"950b80f5",
   506 => x"2d7107b9",
   507 => x"ca0b80f5",
   508 => x"2db9cb0b",
   509 => x"80f52d71",
   510 => x"882b0753",
   511 => x"5f54525a",
   512 => x"56575573",
   513 => x"81abaa2e",
   514 => x"0981068d",
   515 => x"3875519f",
   516 => x"8d2db5a0",
   517 => x"085690a6",
   518 => x"047382d4",
   519 => x"d52e8738",
   520 => x"b1b05190",
   521 => x"e704b5cc",
   522 => x"5275519d",
   523 => x"9b2db5a0",
   524 => x"0855b5a0",
   525 => x"08802e83",
   526 => x"c2388853",
   527 => x"b18c52b6",
   528 => x"9e518e98",
   529 => x"2db5a008",
   530 => x"8938810b",
   531 => x"b9d40c90",
   532 => x"ed048853",
   533 => x"b18052b6",
   534 => x"82518e98",
   535 => x"2db5a008",
   536 => x"802e8a38",
   537 => x"b1d05185",
   538 => x"f32d91c7",
   539 => x"04b9ca0b",
   540 => x"80f52d54",
   541 => x"7380d52e",
   542 => x"09810680",
   543 => x"ca38b9cb",
   544 => x"0b80f52d",
   545 => x"547381aa",
   546 => x"2e098106",
   547 => x"ba38800b",
   548 => x"b5cc0b80",
   549 => x"f52d5654",
   550 => x"7481e92e",
   551 => x"83388154",
   552 => x"7481eb2e",
   553 => x"8c388055",
   554 => x"73752e09",
   555 => x"810682cb",
   556 => x"38b5d70b",
   557 => x"80f52d55",
   558 => x"748d38b5",
   559 => x"d80b80f5",
   560 => x"2d547382",
   561 => x"2e863880",
   562 => x"5593fb04",
   563 => x"b5d90b80",
   564 => x"f52d70b9",
   565 => x"cc0cff05",
   566 => x"b9d00cb5",
   567 => x"da0b80f5",
   568 => x"2db5db0b",
   569 => x"80f52d58",
   570 => x"76057782",
   571 => x"80290570",
   572 => x"b9d80cb5",
   573 => x"dc0b80f5",
   574 => x"2d70b9ec",
   575 => x"0cb9d408",
   576 => x"59575876",
   577 => x"802e81a3",
   578 => x"388853b1",
   579 => x"8c52b69e",
   580 => x"518e982d",
   581 => x"b5a00881",
   582 => x"e238b9cc",
   583 => x"0870842b",
   584 => x"b9f00c70",
   585 => x"b9e80cb5",
   586 => x"f10b80f5",
   587 => x"2db5f00b",
   588 => x"80f52d71",
   589 => x"82802905",
   590 => x"b5f20b80",
   591 => x"f52d7084",
   592 => x"80802912",
   593 => x"b5f30b80",
   594 => x"f52d7081",
   595 => x"800a2912",
   596 => x"70b9f40c",
   597 => x"b9ec0871",
   598 => x"29b9d808",
   599 => x"0570b9dc",
   600 => x"0cb5f90b",
   601 => x"80f52db5",
   602 => x"f80b80f5",
   603 => x"2d718280",
   604 => x"2905b5fa",
   605 => x"0b80f52d",
   606 => x"70848080",
   607 => x"2912b5fb",
   608 => x"0b80f52d",
   609 => x"70982b81",
   610 => x"f00a0672",
   611 => x"0570b9e0",
   612 => x"0cfe117e",
   613 => x"297705b9",
   614 => x"e40c5259",
   615 => x"5243545e",
   616 => x"51525952",
   617 => x"5d575957",
   618 => x"93f904b5",
   619 => x"de0b80f5",
   620 => x"2db5dd0b",
   621 => x"80f52d71",
   622 => x"82802905",
   623 => x"70b9f00c",
   624 => x"70a02983",
   625 => x"ff057089",
   626 => x"2a70b9e8",
   627 => x"0cb5e30b",
   628 => x"80f52db5",
   629 => x"e20b80f5",
   630 => x"2d718280",
   631 => x"290570b9",
   632 => x"f40c7b71",
   633 => x"291e70b9",
   634 => x"e40c7db9",
   635 => x"e00c7305",
   636 => x"b9dc0c55",
   637 => x"5e515155",
   638 => x"55815574",
   639 => x"b5a00c02",
   640 => x"a8050d04",
   641 => x"02ec050d",
   642 => x"7670872c",
   643 => x"7180ff06",
   644 => x"555654b9",
   645 => x"d4088a38",
   646 => x"73882c74",
   647 => x"81ff0654",
   648 => x"55b5cc52",
   649 => x"b9d80815",
   650 => x"519d9b2d",
   651 => x"b5a00854",
   652 => x"b5a00880",
   653 => x"2eb338b9",
   654 => x"d408802e",
   655 => x"98387284",
   656 => x"29b5cc05",
   657 => x"70085253",
   658 => x"9f8d2db5",
   659 => x"a008f00a",
   660 => x"065394e7",
   661 => x"047210b5",
   662 => x"cc057080",
   663 => x"e02d5253",
   664 => x"9fbd2db5",
   665 => x"a0085372",
   666 => x"5473b5a0",
   667 => x"0c029405",
   668 => x"0d0402c8",
   669 => x"050d7f61",
   670 => x"5f5b800b",
   671 => x"b9e008b9",
   672 => x"e408595d",
   673 => x"56b9d408",
   674 => x"762e8a38",
   675 => x"b9cc0884",
   676 => x"2b58959b",
   677 => x"04b9e808",
   678 => x"842b5880",
   679 => x"59787827",
   680 => x"81a93878",
   681 => x"8f06a017",
   682 => x"5754738f",
   683 => x"38b5cc52",
   684 => x"76518117",
   685 => x"579d9b2d",
   686 => x"b5cc5680",
   687 => x"7680f52d",
   688 => x"56547474",
   689 => x"2e833881",
   690 => x"547481e5",
   691 => x"2e80f638",
   692 => x"81707506",
   693 => x"555d7380",
   694 => x"2e80ea38",
   695 => x"8b1680f5",
   696 => x"2d98065a",
   697 => x"7980de38",
   698 => x"8b537d52",
   699 => x"75518e98",
   700 => x"2db5a008",
   701 => x"80cf389c",
   702 => x"1608519f",
   703 => x"8d2db5a0",
   704 => x"08841c0c",
   705 => x"9a1680e0",
   706 => x"2d519fbd",
   707 => x"2db5a008",
   708 => x"b5a00888",
   709 => x"1d0cb5a0",
   710 => x"085555b9",
   711 => x"d408802e",
   712 => x"98389416",
   713 => x"80e02d51",
   714 => x"9fbd2db5",
   715 => x"a008902b",
   716 => x"83fff00a",
   717 => x"06701651",
   718 => x"5473881c",
   719 => x"0c797b0c",
   720 => x"7c549781",
   721 => x"04811959",
   722 => x"959d04b9",
   723 => x"d408802e",
   724 => x"ae387b51",
   725 => x"94842db5",
   726 => x"a008b5a0",
   727 => x"0880ffff",
   728 => x"fff80655",
   729 => x"5c7380ff",
   730 => x"fffff82e",
   731 => x"9238b5a0",
   732 => x"08fe05b9",
   733 => x"cc0829b9",
   734 => x"dc080557",
   735 => x"959b0480",
   736 => x"5473b5a0",
   737 => x"0c02b805",
   738 => x"0d0402f4",
   739 => x"050d7470",
   740 => x"08810571",
   741 => x"0c7008b9",
   742 => x"d0080653",
   743 => x"53718e38",
   744 => x"88130851",
   745 => x"94842db5",
   746 => x"a0088814",
   747 => x"0c810bb5",
   748 => x"a00c028c",
   749 => x"050d0402",
   750 => x"f0050d75",
   751 => x"881108fe",
   752 => x"05b9cc08",
   753 => x"29b9dc08",
   754 => x"117208b9",
   755 => x"d0080605",
   756 => x"79555354",
   757 => x"549d9b2d",
   758 => x"0290050d",
   759 => x"04b9d408",
   760 => x"b5a00c04",
   761 => x"02f4050d",
   762 => x"d45281ff",
   763 => x"720c7108",
   764 => x"5381ff72",
   765 => x"0c72882b",
   766 => x"83fe8006",
   767 => x"72087081",
   768 => x"ff065152",
   769 => x"5381ff72",
   770 => x"0c727107",
   771 => x"882b7208",
   772 => x"7081ff06",
   773 => x"51525381",
   774 => x"ff720c72",
   775 => x"7107882b",
   776 => x"72087081",
   777 => x"ff067207",
   778 => x"b5a00c52",
   779 => x"53028c05",
   780 => x"0d0402f4",
   781 => x"050d7476",
   782 => x"7181ff06",
   783 => x"d40c5353",
   784 => x"b9fc0885",
   785 => x"3871892b",
   786 => x"5271982a",
   787 => x"d40c7190",
   788 => x"2a7081ff",
   789 => x"06d40c51",
   790 => x"71882a70",
   791 => x"81ff06d4",
   792 => x"0c517181",
   793 => x"ff06d40c",
   794 => x"72902a70",
   795 => x"81ff06d4",
   796 => x"0c51d408",
   797 => x"7081ff06",
   798 => x"515182b8",
   799 => x"bf527081",
   800 => x"ff2e0981",
   801 => x"06943881",
   802 => x"ff0bd40c",
   803 => x"d4087081",
   804 => x"ff06ff14",
   805 => x"54515171",
   806 => x"e53870b5",
   807 => x"a00c028c",
   808 => x"050d0402",
   809 => x"fc050d81",
   810 => x"c75181ff",
   811 => x"0bd40cff",
   812 => x"11517080",
   813 => x"25f43802",
   814 => x"84050d04",
   815 => x"02f0050d",
   816 => x"99a32d8f",
   817 => x"cf538052",
   818 => x"87fc80f7",
   819 => x"5198b22d",
   820 => x"b5a00854",
   821 => x"b5a00881",
   822 => x"2e098106",
   823 => x"a33881ff",
   824 => x"0bd40c82",
   825 => x"0a52849c",
   826 => x"80e95198",
   827 => x"b22db5a0",
   828 => x"088b3881",
   829 => x"ff0bd40c",
   830 => x"73539a86",
   831 => x"0499a32d",
   832 => x"ff135372",
   833 => x"c13872b5",
   834 => x"a00c0290",
   835 => x"050d0402",
   836 => x"f4050d81",
   837 => x"ff0bd40c",
   838 => x"93538052",
   839 => x"87fc80c1",
   840 => x"5198b22d",
   841 => x"b5a0088b",
   842 => x"3881ff0b",
   843 => x"d40c8153",
   844 => x"9abc0499",
   845 => x"a32dff13",
   846 => x"5372df38",
   847 => x"72b5a00c",
   848 => x"028c050d",
   849 => x"0402f005",
   850 => x"0d99a32d",
   851 => x"83aa5284",
   852 => x"9c80c851",
   853 => x"98b22db5",
   854 => x"a008812e",
   855 => x"09810692",
   856 => x"3897e42d",
   857 => x"b5a00883",
   858 => x"ffff0653",
   859 => x"7283aa2e",
   860 => x"97389a8f",
   861 => x"2d9b8304",
   862 => x"81549bf2",
   863 => x"04b1f051",
   864 => x"85f32d80",
   865 => x"549bf204",
   866 => x"81ff0bd4",
   867 => x"0cb15399",
   868 => x"bc2db5a0",
   869 => x"08802e80",
   870 => x"ca388052",
   871 => x"87fc80fa",
   872 => x"5198b22d",
   873 => x"b5a008b1",
   874 => x"3881ff0b",
   875 => x"d40cd408",
   876 => x"5381ff0b",
   877 => x"d40c81ff",
   878 => x"0bd40c81",
   879 => x"ff0bd40c",
   880 => x"81ff0bd4",
   881 => x"0c72862a",
   882 => x"708106b5",
   883 => x"a0085651",
   884 => x"5372802e",
   885 => x"9d389af8",
   886 => x"04b5a008",
   887 => x"52b28c51",
   888 => x"a0b82d72",
   889 => x"822eff95",
   890 => x"38ff1353",
   891 => x"72ffa038",
   892 => x"725473b5",
   893 => x"a00c0290",
   894 => x"050d0402",
   895 => x"f4050d81",
   896 => x"0bb9fc0c",
   897 => x"d008708f",
   898 => x"2a708106",
   899 => x"51515372",
   900 => x"f33872d0",
   901 => x"0c99a32d",
   902 => x"b2985185",
   903 => x"f32dd008",
   904 => x"708f2a70",
   905 => x"81065151",
   906 => x"5372f338",
   907 => x"810bd00c",
   908 => x"80e35380",
   909 => x"5284d480",
   910 => x"c05198b2",
   911 => x"2db5a008",
   912 => x"812e9a38",
   913 => x"72822e09",
   914 => x"81068c38",
   915 => x"b2b45185",
   916 => x"f32d8053",
   917 => x"9d9204ff",
   918 => x"135372d7",
   919 => x"389ac52d",
   920 => x"b5a008b9",
   921 => x"fc0cb5a0",
   922 => x"088b3881",
   923 => x"5287fc80",
   924 => x"d05198b2",
   925 => x"2d81ff0b",
   926 => x"d40cd008",
   927 => x"708f2a70",
   928 => x"81065151",
   929 => x"5372f338",
   930 => x"72d00c81",
   931 => x"ff0bd40c",
   932 => x"815372b5",
   933 => x"a00c028c",
   934 => x"050d0402",
   935 => x"e0050d79",
   936 => x"7b575780",
   937 => x"5881ff0b",
   938 => x"d40cd008",
   939 => x"708f2a70",
   940 => x"81065151",
   941 => x"5473f338",
   942 => x"82810bd0",
   943 => x"0c81ff0b",
   944 => x"d40c7652",
   945 => x"87fc80d1",
   946 => x"5198b22d",
   947 => x"80dbc6df",
   948 => x"55b5a008",
   949 => x"802e9038",
   950 => x"b5a00853",
   951 => x"7652b2cc",
   952 => x"51a0b82d",
   953 => x"9eb50481",
   954 => x"ff0bd40c",
   955 => x"d4087081",
   956 => x"ff065154",
   957 => x"7381fe2e",
   958 => x"0981069d",
   959 => x"3880ff54",
   960 => x"97e42db5",
   961 => x"a0087670",
   962 => x"8405580c",
   963 => x"ff145473",
   964 => x"8025ed38",
   965 => x"81589e9f",
   966 => x"04ff1555",
   967 => x"74c93881",
   968 => x"ff0bd40c",
   969 => x"d008708f",
   970 => x"2a708106",
   971 => x"51515473",
   972 => x"f33873d0",
   973 => x"0c77b5a0",
   974 => x"0c02a005",
   975 => x"0d04b9fc",
   976 => x"08b5a00c",
   977 => x"0402e805",
   978 => x"0d807857",
   979 => x"55757084",
   980 => x"05570853",
   981 => x"80547298",
   982 => x"2a73882b",
   983 => x"54527180",
   984 => x"2ea238c0",
   985 => x"0870882a",
   986 => x"70810651",
   987 => x"51517080",
   988 => x"2ef13871",
   989 => x"c00c8115",
   990 => x"81155555",
   991 => x"837425d6",
   992 => x"3871ca38",
   993 => x"74b5a00c",
   994 => x"0298050d",
   995 => x"0402f405",
   996 => x"0d747088",
   997 => x"2a83fe80",
   998 => x"06707298",
   999 => x"2a077288",
  1000 => x"2b87fc80",
  1001 => x"80067398",
  1002 => x"2b81f00a",
  1003 => x"06717307",
  1004 => x"07b5a00c",
  1005 => x"56515351",
  1006 => x"028c050d",
  1007 => x"0402f805",
  1008 => x"0d028e05",
  1009 => x"80f52d74",
  1010 => x"882b0770",
  1011 => x"83ffff06",
  1012 => x"b5a00c51",
  1013 => x"0288050d",
  1014 => x"0402ec05",
  1015 => x"0d765380",
  1016 => x"55727525",
  1017 => x"8b38ad51",
  1018 => x"82ee2d72",
  1019 => x"09810553",
  1020 => x"72802eb5",
  1021 => x"38875472",
  1022 => x"9c2a7384",
  1023 => x"2b545271",
  1024 => x"802e8338",
  1025 => x"81558972",
  1026 => x"258738b7",
  1027 => x"1252a094",
  1028 => x"04b01252",
  1029 => x"74802e86",
  1030 => x"38715182",
  1031 => x"ee2dff14",
  1032 => x"54738025",
  1033 => x"d238a0ae",
  1034 => x"04b05182",
  1035 => x"ee2d800b",
  1036 => x"b5a00c02",
  1037 => x"94050d04",
  1038 => x"02c0050d",
  1039 => x"0280c405",
  1040 => x"57807078",
  1041 => x"7084055a",
  1042 => x"0872415f",
  1043 => x"5d587c70",
  1044 => x"84055e08",
  1045 => x"5a805b79",
  1046 => x"982a7a88",
  1047 => x"2b5b5675",
  1048 => x"8638775f",
  1049 => x"a2b0047d",
  1050 => x"802e81a2",
  1051 => x"38805e75",
  1052 => x"80e42e8a",
  1053 => x"387580f8",
  1054 => x"2e098106",
  1055 => x"89387684",
  1056 => x"1871085e",
  1057 => x"58547580",
  1058 => x"e42e9f38",
  1059 => x"7580e426",
  1060 => x"8a387580",
  1061 => x"e32ebe38",
  1062 => x"a1e00475",
  1063 => x"80f32ea3",
  1064 => x"387580f8",
  1065 => x"2e8938a1",
  1066 => x"e0048a53",
  1067 => x"a1b10490",
  1068 => x"53ba8052",
  1069 => x"7b519fd9",
  1070 => x"2db5a008",
  1071 => x"ba805a55",
  1072 => x"a1f00476",
  1073 => x"84187108",
  1074 => x"70545b58",
  1075 => x"549ec52d",
  1076 => x"8055a1f0",
  1077 => x"04768418",
  1078 => x"71085858",
  1079 => x"54a29b04",
  1080 => x"a55182ee",
  1081 => x"2d755182",
  1082 => x"ee2d8218",
  1083 => x"58a2a304",
  1084 => x"74ff1656",
  1085 => x"54807425",
  1086 => x"aa387870",
  1087 => x"81055a80",
  1088 => x"f52d7052",
  1089 => x"5682ee2d",
  1090 => x"811858a1",
  1091 => x"f00475a5",
  1092 => x"2e098106",
  1093 => x"8638815e",
  1094 => x"a2a30475",
  1095 => x"5182ee2d",
  1096 => x"81185881",
  1097 => x"1b5b837b",
  1098 => x"25feac38",
  1099 => x"75fe9f38",
  1100 => x"7eb5a00c",
  1101 => x"0280c005",
  1102 => x"0d0402fc",
  1103 => x"050d7251",
  1104 => x"80710c80",
  1105 => x"0b84120c",
  1106 => x"0284050d",
  1107 => x"0402f005",
  1108 => x"0d757008",
  1109 => x"84120853",
  1110 => x"5353ff54",
  1111 => x"71712ea8",
  1112 => x"38a7be2d",
  1113 => x"84130870",
  1114 => x"84291488",
  1115 => x"11700870",
  1116 => x"81ff0684",
  1117 => x"18088111",
  1118 => x"8706841a",
  1119 => x"0c535155",
  1120 => x"515151a7",
  1121 => x"b82d7154",
  1122 => x"73b5a00c",
  1123 => x"0290050d",
  1124 => x"0402f405",
  1125 => x"0d745384",
  1126 => x"13088111",
  1127 => x"87067408",
  1128 => x"54515171",
  1129 => x"712ef038",
  1130 => x"a7be2d84",
  1131 => x"13087084",
  1132 => x"29148811",
  1133 => x"78710c51",
  1134 => x"51518413",
  1135 => x"08811187",
  1136 => x"0684150c",
  1137 => x"51a7b82d",
  1138 => x"028c050d",
  1139 => x"0402f405",
  1140 => x"0da7be2d",
  1141 => x"e008e408",
  1142 => x"718b2a70",
  1143 => x"81065153",
  1144 => x"54527080",
  1145 => x"2e9d38ba",
  1146 => x"c0087084",
  1147 => x"29bac805",
  1148 => x"7381ff06",
  1149 => x"710c5151",
  1150 => x"bac00881",
  1151 => x"118706ba",
  1152 => x"c00c5172",
  1153 => x"8b2a7081",
  1154 => x"06515170",
  1155 => x"802eb238",
  1156 => x"bae80870",
  1157 => x"8429baf0",
  1158 => x"057481ff",
  1159 => x"06710c51",
  1160 => x"51bae808",
  1161 => x"81118706",
  1162 => x"bae80c51",
  1163 => x"bae808ba",
  1164 => x"ec085252",
  1165 => x"71712e09",
  1166 => x"81068638",
  1167 => x"810bbbb8",
  1168 => x"0c728a2a",
  1169 => x"70810651",
  1170 => x"5170802e",
  1171 => x"a838bb90",
  1172 => x"08bb9408",
  1173 => x"52527171",
  1174 => x"2e9b38bb",
  1175 => x"90087084",
  1176 => x"29bb9805",
  1177 => x"7008e40c",
  1178 => x"5151bb90",
  1179 => x"08811187",
  1180 => x"06bb900c",
  1181 => x"51800bbb",
  1182 => x"bc0ca7b1",
  1183 => x"2da7b82d",
  1184 => x"028c050d",
  1185 => x"0402fc05",
  1186 => x"0da7be2d",
  1187 => x"810bbbbc",
  1188 => x"0ca7b82d",
  1189 => x"bbbc0851",
  1190 => x"70fa3802",
  1191 => x"84050d04",
  1192 => x"02fc050d",
  1193 => x"800bbbb8",
  1194 => x"0cbac051",
  1195 => x"a2ba2da3",
  1196 => x"cd51a7ad",
  1197 => x"2da6d72d",
  1198 => x"0284050d",
  1199 => x"0402f405",
  1200 => x"0da6bf04",
  1201 => x"b5a00881",
  1202 => x"f02e0981",
  1203 => x"06893881",
  1204 => x"0bb5940c",
  1205 => x"a6bf04b5",
  1206 => x"a00881e0",
  1207 => x"2e098106",
  1208 => x"8938810b",
  1209 => x"b5980ca6",
  1210 => x"bf04b5a0",
  1211 => x"0852b598",
  1212 => x"08802e88",
  1213 => x"38b5a008",
  1214 => x"81800552",
  1215 => x"71842c72",
  1216 => x"8f065353",
  1217 => x"b5940880",
  1218 => x"2e993872",
  1219 => x"8429b4d4",
  1220 => x"05721381",
  1221 => x"712b7009",
  1222 => x"73080673",
  1223 => x"0c515353",
  1224 => x"a6b50472",
  1225 => x"8429b4d4",
  1226 => x"05721383",
  1227 => x"712b7208",
  1228 => x"07720c53",
  1229 => x"53800bb5",
  1230 => x"980c800b",
  1231 => x"b5940cba",
  1232 => x"c051a2cd",
  1233 => x"2db5a008",
  1234 => x"ff24fef8",
  1235 => x"38800bb5",
  1236 => x"a00c028c",
  1237 => x"050d0402",
  1238 => x"f8050db4",
  1239 => x"d4528f51",
  1240 => x"80727084",
  1241 => x"05540cff",
  1242 => x"11517080",
  1243 => x"25f23802",
  1244 => x"88050d04",
  1245 => x"02f0050d",
  1246 => x"7551a7be",
  1247 => x"2d70822c",
  1248 => x"fc06b4d4",
  1249 => x"1172109e",
  1250 => x"06710870",
  1251 => x"722a7083",
  1252 => x"0682742b",
  1253 => x"70097406",
  1254 => x"760c5451",
  1255 => x"56575351",
  1256 => x"53a7b82d",
  1257 => x"71b5a00c",
  1258 => x"0290050d",
  1259 => x"0471980c",
  1260 => x"04ffb008",
  1261 => x"b5a00c04",
  1262 => x"810bffb0",
  1263 => x"0c04800b",
  1264 => x"ffb00c04",
  1265 => x"02fc050d",
  1266 => x"800bb59c",
  1267 => x"0c805184",
  1268 => x"e52d0284",
  1269 => x"050d0402",
  1270 => x"f0050dbb",
  1271 => x"c4085481",
  1272 => x"f72d800b",
  1273 => x"bbc80c73",
  1274 => x"08802e80",
  1275 => x"eb38820b",
  1276 => x"b5b40cbb",
  1277 => x"c8088f06",
  1278 => x"b5b00c73",
  1279 => x"08527181",
  1280 => x"2ea43871",
  1281 => x"832e0981",
  1282 => x"06b93888",
  1283 => x"1480f52d",
  1284 => x"841508b2",
  1285 => x"ec535452",
  1286 => x"85f32d71",
  1287 => x"84291370",
  1288 => x"085252a8",
  1289 => x"c704bbc0",
  1290 => x"08881508",
  1291 => x"2c708106",
  1292 => x"51527180",
  1293 => x"2e8738b2",
  1294 => x"f051a8c0",
  1295 => x"04b2f451",
  1296 => x"85f32d84",
  1297 => x"14085185",
  1298 => x"f32dbbc8",
  1299 => x"088105bb",
  1300 => x"c80c8c14",
  1301 => x"54a7e704",
  1302 => x"0290050d",
  1303 => x"0471bbc4",
  1304 => x"0ca7d72d",
  1305 => x"bbc808ff",
  1306 => x"05bbcc0c",
  1307 => x"0402f005",
  1308 => x"0d8751a6",
  1309 => x"f42db5a0",
  1310 => x"08812a70",
  1311 => x"81065152",
  1312 => x"71802ea0",
  1313 => x"38a98b04",
  1314 => x"a5bd2d87",
  1315 => x"51a6f42d",
  1316 => x"b5a008f4",
  1317 => x"38b59c08",
  1318 => x"813270b5",
  1319 => x"9c0c7052",
  1320 => x"5284e52d",
  1321 => x"b59c0896",
  1322 => x"3880da51",
  1323 => x"a6f42d81",
  1324 => x"f551a6f4",
  1325 => x"2d81f251",
  1326 => x"a6f42dab",
  1327 => x"db0481f5",
  1328 => x"51a6f42d",
  1329 => x"b5a00881",
  1330 => x"2a708106",
  1331 => x"51527180",
  1332 => x"2e8f38bb",
  1333 => x"cc085271",
  1334 => x"802e8638",
  1335 => x"ff12bbcc",
  1336 => x"0c81f251",
  1337 => x"a6f42db5",
  1338 => x"a008812a",
  1339 => x"70810651",
  1340 => x"5271802e",
  1341 => x"9538bbc8",
  1342 => x"08ff05bb",
  1343 => x"cc085452",
  1344 => x"72722586",
  1345 => x"388113bb",
  1346 => x"cc0c80da",
  1347 => x"51a6f42d",
  1348 => x"b5a00881",
  1349 => x"2a708106",
  1350 => x"51527180",
  1351 => x"2e80fb38",
  1352 => x"bbc408bb",
  1353 => x"cc085553",
  1354 => x"73802e8a",
  1355 => x"388c13ff",
  1356 => x"155553aa",
  1357 => x"a8047208",
  1358 => x"5271822e",
  1359 => x"a6387182",
  1360 => x"26893871",
  1361 => x"812ea538",
  1362 => x"ab9a0471",
  1363 => x"832ead38",
  1364 => x"71842e09",
  1365 => x"810680c2",
  1366 => x"38881308",
  1367 => x"51a8dd2d",
  1368 => x"ab9a0488",
  1369 => x"13085271",
  1370 => x"2dab9a04",
  1371 => x"810b8814",
  1372 => x"082bbbc0",
  1373 => x"0832bbc0",
  1374 => x"0cab9704",
  1375 => x"881380f5",
  1376 => x"2d81058b",
  1377 => x"1480f52d",
  1378 => x"53547174",
  1379 => x"24833880",
  1380 => x"54738814",
  1381 => x"81b72da7",
  1382 => x"d72d8054",
  1383 => x"800bb5b4",
  1384 => x"0c738f06",
  1385 => x"b5b00ca0",
  1386 => x"5273bbcc",
  1387 => x"082e0981",
  1388 => x"069838bb",
  1389 => x"c808ff05",
  1390 => x"74327009",
  1391 => x"81057072",
  1392 => x"079f2a91",
  1393 => x"71315151",
  1394 => x"53537151",
  1395 => x"82ee2d81",
  1396 => x"14548e74",
  1397 => x"25c638b5",
  1398 => x"9c085271",
  1399 => x"b5a00c02",
  1400 => x"90050d04",
  1401 => x"00ffffff",
  1402 => x"ff00ffff",
  1403 => x"ffff00ff",
  1404 => x"ffffff00",
  1405 => x"52657365",
  1406 => x"74000000",
  1407 => x"4f707469",
  1408 => x"6f6e7320",
  1409 => x"10000000",
  1410 => x"54757262",
  1411 => x"6f202831",
  1412 => x"302e3734",
  1413 => x"4d487a29",
  1414 => x"00000000",
  1415 => x"4d6f7573",
  1416 => x"6520656d",
  1417 => x"756c6174",
  1418 => x"696f6e00",
  1419 => x"45786974",
  1420 => x"00000000",
  1421 => x"53442043",
  1422 => x"61726400",
  1423 => x"4a617061",
  1424 => x"6e657365",
  1425 => x"206b6579",
  1426 => x"626f6172",
  1427 => x"64206c61",
  1428 => x"796f7574",
  1429 => x"00000000",
  1430 => x"4261636b",
  1431 => x"00000000",
  1432 => x"32303438",
  1433 => x"4c422052",
  1434 => x"414d0000",
  1435 => x"34303936",
  1436 => x"4b422052",
  1437 => x"414d0000",
  1438 => x"536c323a",
  1439 => x"204e6f6e",
  1440 => x"65000000",
  1441 => x"536c323a",
  1442 => x"20455345",
  1443 => x"2d534343",
  1444 => x"20314d42",
  1445 => x"2f534343",
  1446 => x"2d490000",
  1447 => x"536c323a",
  1448 => x"20455345",
  1449 => x"2d52414d",
  1450 => x"20314d42",
  1451 => x"2f415343",
  1452 => x"49493800",
  1453 => x"536c323a",
  1454 => x"20455345",
  1455 => x"2d52414d",
  1456 => x"20314d42",
  1457 => x"2f415343",
  1458 => x"49493136",
  1459 => x"00000000",
  1460 => x"536c313a",
  1461 => x"204e6f6e",
  1462 => x"65000000",
  1463 => x"536c313a",
  1464 => x"20455345",
  1465 => x"2d534343",
  1466 => x"20314d42",
  1467 => x"2f534343",
  1468 => x"2d490000",
  1469 => x"536c313a",
  1470 => x"204d6567",
  1471 => x"6152414d",
  1472 => x"00000000",
  1473 => x"56474120",
  1474 => x"2d203331",
  1475 => x"4b487a2c",
  1476 => x"20363048",
  1477 => x"7a000000",
  1478 => x"56474120",
  1479 => x"2d203331",
  1480 => x"4b487a2c",
  1481 => x"20353048",
  1482 => x"7a000000",
  1483 => x"5456202d",
  1484 => x"20343830",
  1485 => x"692c2036",
  1486 => x"30487a00",
  1487 => x"496e6974",
  1488 => x"69616c69",
  1489 => x"7a696e67",
  1490 => x"20534420",
  1491 => x"63617264",
  1492 => x"0a000000",
  1493 => x"53444843",
  1494 => x"20636172",
  1495 => x"64206465",
  1496 => x"74656374",
  1497 => x"65642062",
  1498 => x"7574206e",
  1499 => x"6f740a73",
  1500 => x"7570706f",
  1501 => x"72746564",
  1502 => x"3b206469",
  1503 => x"7361626c",
  1504 => x"696e6720",
  1505 => x"53442063",
  1506 => x"6172640a",
  1507 => x"10204f4b",
  1508 => x"0a000000",
  1509 => x"46617433",
  1510 => x"32206669",
  1511 => x"6c657379",
  1512 => x"7374656d",
  1513 => x"20646574",
  1514 => x"65637465",
  1515 => x"64206275",
  1516 => x"740a6e6f",
  1517 => x"74207375",
  1518 => x"70706f72",
  1519 => x"7465643b",
  1520 => x"20646973",
  1521 => x"61626c69",
  1522 => x"6e672053",
  1523 => x"44206361",
  1524 => x"72640a10",
  1525 => x"204f4b0a",
  1526 => x"00000000",
  1527 => x"54727969",
  1528 => x"6e67204d",
  1529 => x"53583342",
  1530 => x"494f532e",
  1531 => x"5359532e",
  1532 => x"2e2e0a00",
  1533 => x"4d535833",
  1534 => x"42494f53",
  1535 => x"53595300",
  1536 => x"54727969",
  1537 => x"6e672042",
  1538 => x"494f535f",
  1539 => x"4d32502e",
  1540 => x"524f4d2e",
  1541 => x"2e2e0a00",
  1542 => x"42494f53",
  1543 => x"5f4d3250",
  1544 => x"524f4d00",
  1545 => x"4f70656e",
  1546 => x"65642042",
  1547 => x"494f532c",
  1548 => x"206c6f61",
  1549 => x"64696e67",
  1550 => x"2e2e2e0a",
  1551 => x"00000000",
  1552 => x"52656164",
  1553 => x"20626c6f",
  1554 => x"636b2066",
  1555 => x"61696c65",
  1556 => x"640a0000",
  1557 => x"4c6f6164",
  1558 => x"696e6720",
  1559 => x"42494f53",
  1560 => x"20666169",
  1561 => x"6c65640a",
  1562 => x"00000000",
  1563 => x"52656164",
  1564 => x"206f6620",
  1565 => x"4d425220",
  1566 => x"6661696c",
  1567 => x"65640a00",
  1568 => x"46415431",
  1569 => x"36202020",
  1570 => x"00000000",
  1571 => x"46415433",
  1572 => x"32202020",
  1573 => x"00000000",
  1574 => x"25642070",
  1575 => x"61727469",
  1576 => x"74696f6e",
  1577 => x"7320666f",
  1578 => x"756e640a",
  1579 => x"00000000",
  1580 => x"4e6f2070",
  1581 => x"61727469",
  1582 => x"74696f6e",
  1583 => x"20736967",
  1584 => x"6e617475",
  1585 => x"72652066",
  1586 => x"6f756e64",
  1587 => x"0a000000",
  1588 => x"556e7375",
  1589 => x"70706f72",
  1590 => x"74656420",
  1591 => x"70617274",
  1592 => x"6974696f",
  1593 => x"6e207479",
  1594 => x"7065210a",
  1595 => x"00000000",
  1596 => x"53444843",
  1597 => x"20496e69",
  1598 => x"7469616c",
  1599 => x"697a6174",
  1600 => x"696f6e20",
  1601 => x"6572726f",
  1602 => x"72210a00",
  1603 => x"434d4435",
  1604 => x"38202564",
  1605 => x"0a202000",
  1606 => x"496e6974",
  1607 => x"69616c69",
  1608 => x"7a696e67",
  1609 => x"20534420",
  1610 => x"63617264",
  1611 => x"2e2e2e0a",
  1612 => x"00000000",
  1613 => x"53442063",
  1614 => x"61726420",
  1615 => x"72657365",
  1616 => x"74206661",
  1617 => x"696c6564",
  1618 => x"210a0000",
  1619 => x"52656164",
  1620 => x"20636f6d",
  1621 => x"6d616e64",
  1622 => x"20666169",
  1623 => x"6c656420",
  1624 => x"61742025",
  1625 => x"64202825",
  1626 => x"64290a00",
  1627 => x"16200000",
  1628 => x"14200000",
  1629 => x"15200000",
  1630 => x"00000002",
  1631 => x"00000002",
  1632 => x"000015f4",
  1633 => x"00000540",
  1634 => x"00000004",
  1635 => x"000015fc",
  1636 => x"000019c4",
  1637 => x"00000001",
  1638 => x"00001608",
  1639 => x"00000007",
  1640 => x"00000001",
  1641 => x"0000161c",
  1642 => x"0000000a",
  1643 => x"00000002",
  1644 => x"0000162c",
  1645 => x"000013c4",
  1646 => x"00000000",
  1647 => x"00000000",
  1648 => x"00000000",
  1649 => x"00000003",
  1650 => x"00001a48",
  1651 => x"00000003",
  1652 => x"00000001",
  1653 => x"00001634",
  1654 => x"00000002",
  1655 => x"00000003",
  1656 => x"00001a3c",
  1657 => x"00000003",
  1658 => x"00000003",
  1659 => x"00001a2c",
  1660 => x"00000004",
  1661 => x"00000001",
  1662 => x"0000163c",
  1663 => x"00000006",
  1664 => x"00000003",
  1665 => x"00001a24",
  1666 => x"00000002",
  1667 => x"00000004",
  1668 => x"00001658",
  1669 => x"0000197c",
  1670 => x"00000000",
  1671 => x"00000000",
  1672 => x"00000000",
  1673 => x"00001660",
  1674 => x"0000166c",
  1675 => x"00001678",
  1676 => x"00001684",
  1677 => x"0000169c",
  1678 => x"000016b4",
  1679 => x"000016d0",
  1680 => x"000016dc",
  1681 => x"000016f4",
  1682 => x"00001704",
  1683 => x"00001718",
  1684 => x"0000172c",
  1685 => x"00000000",
  1686 => x"00000000",
  1687 => x"00000000",
  1688 => x"00000000",
  1689 => x"00000000",
  1690 => x"00000000",
  1691 => x"00000000",
  1692 => x"00000000",
  1693 => x"00000000",
  1694 => x"00000000",
  1695 => x"00000000",
  1696 => x"00000000",
  1697 => x"00000000",
  1698 => x"00000000",
  1699 => x"00000000",
  1700 => x"00000000",
  1701 => x"00000000",
  1702 => x"00000000",
  1703 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

