-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"000b0b0b",
     4 => x"0b8c04ff",
     5 => x"0d800404",
     6 => x"00000017",
     7 => x"00000000",
     8 => x"0b0b0bba",
     9 => x"ac080b0b",
    10 => x"0bbab008",
    11 => x"0b0b0bba",
    12 => x"b4080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"bab40c0b",
    16 => x"0b0bbab0",
    17 => x"0c0b0b0b",
    18 => x"baac0c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0bb098",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"baac70bf",
    57 => x"e4278b38",
    58 => x"80717084",
    59 => x"05530c81",
    60 => x"e2048c51",
    61 => x"8dec0402",
    62 => x"fc050df8",
    63 => x"80518f0b",
    64 => x"babc0c9f",
    65 => x"0bbac00c",
    66 => x"a0717081",
    67 => x"055334ba",
    68 => x"c008ff05",
    69 => x"bac00cba",
    70 => x"c0088025",
    71 => x"eb38babc",
    72 => x"08ff05ba",
    73 => x"bc0cbabc",
    74 => x"088025d7",
    75 => x"38028405",
    76 => x"0d0402f0",
    77 => x"050df880",
    78 => x"53f8a054",
    79 => x"83bf5273",
    80 => x"70810555",
    81 => x"33517073",
    82 => x"70810555",
    83 => x"34ff1252",
    84 => x"718025eb",
    85 => x"38fbc053",
    86 => x"9f52a073",
    87 => x"70810555",
    88 => x"34ff1252",
    89 => x"718025f2",
    90 => x"38029005",
    91 => x"0d0402f4",
    92 => x"050d7453",
    93 => x"8e0bbabc",
    94 => x"08258f38",
    95 => x"82b22dba",
    96 => x"bc08ff05",
    97 => x"babc0c82",
    98 => x"f404babc",
    99 => x"08bac008",
   100 => x"5351728a",
   101 => x"2e098106",
   102 => x"b7387151",
   103 => x"719f24a0",
   104 => x"38babc08",
   105 => x"a02911f8",
   106 => x"80115151",
   107 => x"a07134ba",
   108 => x"c0088105",
   109 => x"bac00cba",
   110 => x"c008519f",
   111 => x"7125e238",
   112 => x"800bbac0",
   113 => x"0cbabc08",
   114 => x"8105babc",
   115 => x"0c83e404",
   116 => x"70a02912",
   117 => x"f8801151",
   118 => x"51727134",
   119 => x"bac00881",
   120 => x"05bac00c",
   121 => x"bac008a0",
   122 => x"2e098106",
   123 => x"8e38800b",
   124 => x"bac00cba",
   125 => x"bc088105",
   126 => x"babc0c02",
   127 => x"8c050d04",
   128 => x"02e8050d",
   129 => x"77795656",
   130 => x"880bfc16",
   131 => x"77712c8f",
   132 => x"06545254",
   133 => x"80537272",
   134 => x"25953871",
   135 => x"53fbe014",
   136 => x"51877134",
   137 => x"8114ff14",
   138 => x"545472f1",
   139 => x"387153f9",
   140 => x"1576712c",
   141 => x"87065351",
   142 => x"71802e8b",
   143 => x"38fbe014",
   144 => x"51717134",
   145 => x"81145472",
   146 => x"8e249538",
   147 => x"8f733153",
   148 => x"fbe01451",
   149 => x"a0713481",
   150 => x"14ff1454",
   151 => x"5472f138",
   152 => x"0298050d",
   153 => x"0402ec05",
   154 => x"0d800bba",
   155 => x"c40cf68c",
   156 => x"08f69008",
   157 => x"71882c56",
   158 => x"5481ff06",
   159 => x"52737225",
   160 => x"88387154",
   161 => x"820bbac4",
   162 => x"0c72882c",
   163 => x"7381ff06",
   164 => x"54557473",
   165 => x"258b3872",
   166 => x"bac40884",
   167 => x"07bac40c",
   168 => x"5573842b",
   169 => x"86a07125",
   170 => x"83713170",
   171 => x"0b0b0bb6",
   172 => x"e40c8171",
   173 => x"2bff05f6",
   174 => x"880cfecc",
   175 => x"13ff122c",
   176 => x"788829ff",
   177 => x"94057081",
   178 => x"2cbac408",
   179 => x"52585255",
   180 => x"51525476",
   181 => x"802e8538",
   182 => x"70810751",
   183 => x"70f6940c",
   184 => x"71098105",
   185 => x"f6800c72",
   186 => x"098105f6",
   187 => x"840c0294",
   188 => x"050d0402",
   189 => x"f4050d74",
   190 => x"53727081",
   191 => x"055480f5",
   192 => x"2d527180",
   193 => x"2e893871",
   194 => x"5182ee2d",
   195 => x"85f90402",
   196 => x"8c050d04",
   197 => x"02f8050d",
   198 => x"a7ad2d80",
   199 => x"da51a8e4",
   200 => x"2dbaac08",
   201 => x"812a7081",
   202 => x"06515271",
   203 => x"802ee938",
   204 => x"0288050d",
   205 => x"0402f405",
   206 => x"0dbfd408",
   207 => x"99c406b9",
   208 => x"880b80f5",
   209 => x"2d525270",
   210 => x"802e8638",
   211 => x"71848007",
   212 => x"52b8c00b",
   213 => x"80f52d72",
   214 => x"07b8e40b",
   215 => x"80f52d70",
   216 => x"812a7081",
   217 => x"06515354",
   218 => x"5270802e",
   219 => x"86387182",
   220 => x"80075272",
   221 => x"81065170",
   222 => x"802e8538",
   223 => x"71880752",
   224 => x"b8f00b80",
   225 => x"f52d7084",
   226 => x"2b730781",
   227 => x"8432baac",
   228 => x"0c51028c",
   229 => x"050d0402",
   230 => x"f4050d74",
   231 => x"70818432",
   232 => x"bfd40c70",
   233 => x"83065253",
   234 => x"70b8b80b",
   235 => x"880581b7",
   236 => x"2d72892a",
   237 => x"70810651",
   238 => x"5170b988",
   239 => x"0b81b72d",
   240 => x"72832a81",
   241 => x"0673882a",
   242 => x"70810651",
   243 => x"52527080",
   244 => x"2e853871",
   245 => x"82075271",
   246 => x"b8e40b81",
   247 => x"b72d7284",
   248 => x"2c708306",
   249 => x"515170b8",
   250 => x"f00b81b7",
   251 => x"2d70baac",
   252 => x"0c028c05",
   253 => x"0d0402f4",
   254 => x"050db7f0",
   255 => x"0b881180",
   256 => x"f52d8c12",
   257 => x"881180f5",
   258 => x"2d70842b",
   259 => x"73078c13",
   260 => x"881180f5",
   261 => x"2d70882b",
   262 => x"73079413",
   263 => x"80f52d70",
   264 => x"8c2b7207",
   265 => x"baac0c53",
   266 => x"53535353",
   267 => x"56525351",
   268 => x"028c050d",
   269 => x"04b7a00b",
   270 => x"80f52dba",
   271 => x"ac0c0402",
   272 => x"f4050d74",
   273 => x"b7f07187",
   274 => x"06555351",
   275 => x"72881381",
   276 => x"b72d8c12",
   277 => x"71842c70",
   278 => x"87065552",
   279 => x"52728813",
   280 => x"81b72d8c",
   281 => x"1271842c",
   282 => x"70870655",
   283 => x"52527288",
   284 => x"1381b72d",
   285 => x"70842c70",
   286 => x"87065151",
   287 => x"70941381",
   288 => x"b72d028c",
   289 => x"050d0402",
   290 => x"fc050d02",
   291 => x"8b0580f5",
   292 => x"2db7a00b",
   293 => x"81b72d70",
   294 => x"baac0c02",
   295 => x"84050d04",
   296 => x"02d4050d",
   297 => x"7cb3e452",
   298 => x"5585f32d",
   299 => x"9ed52dba",
   300 => x"ac08802e",
   301 => x"83bd3886",
   302 => x"b52dbaac",
   303 => x"0853919e",
   304 => x"2dbaac08",
   305 => x"54baac08",
   306 => x"802e83a9",
   307 => x"38a2d82d",
   308 => x"baac0880",
   309 => x"2e8738b3",
   310 => x"fc5189ea",
   311 => x"049ac12d",
   312 => x"baac0880",
   313 => x"2ea238b4",
   314 => x"905185f3",
   315 => x"2db4a851",
   316 => x"85f32d86",
   317 => x"942d7284",
   318 => x"0753810b",
   319 => x"fec40c72",
   320 => x"fec00c72",
   321 => x"5187972d",
   322 => x"840bfec4",
   323 => x"0cb4c452",
   324 => x"bacc5197",
   325 => x"b02dbaac",
   326 => x"08802e80",
   327 => x"ec387482",
   328 => x"2e098106",
   329 => x"b83872ba",
   330 => x"d80c87f6",
   331 => x"2dbaac08",
   332 => x"badc0c88",
   333 => x"b52dbaac",
   334 => x"08bae00c",
   335 => x"bae45480",
   336 => x"fc538074",
   337 => x"70840556",
   338 => x"0cff1353",
   339 => x"728025f2",
   340 => x"38bad852",
   341 => x"bacc519a",
   342 => x"9b2d8b89",
   343 => x"0474812e",
   344 => x"098106a5",
   345 => x"38bad852",
   346 => x"bacc5199",
   347 => x"f52dbad8",
   348 => x"08badc08",
   349 => x"525388bf",
   350 => x"2dbae008",
   351 => x"5189872d",
   352 => x"72fec00c",
   353 => x"72518797",
   354 => x"2d7d8938",
   355 => x"810bfec8",
   356 => x"0c8ce904",
   357 => x"b4d05185",
   358 => x"f32db4e8",
   359 => x"52bacc51",
   360 => x"97b02dba",
   361 => x"ac089838",
   362 => x"b4f45185",
   363 => x"f32db58c",
   364 => x"52bacc51",
   365 => x"97b02dba",
   366 => x"ac08802e",
   367 => x"81b538b5",
   368 => x"985185f3",
   369 => x"2dbad008",
   370 => x"57807759",
   371 => x"5a767a2e",
   372 => x"8b38811a",
   373 => x"78812a59",
   374 => x"5a77f738",
   375 => x"f71a5a80",
   376 => x"0bfec80c",
   377 => x"80772581",
   378 => x"80387952",
   379 => x"77518480",
   380 => x"2dbad852",
   381 => x"bacc5199",
   382 => x"f52dbaac",
   383 => x"0853baac",
   384 => x"08802e80",
   385 => x"c938bad8",
   386 => x"5b80598c",
   387 => x"bb047a70",
   388 => x"84055c08",
   389 => x"7081ff06",
   390 => x"71882c70",
   391 => x"81ff0673",
   392 => x"902c7081",
   393 => x"ff067598",
   394 => x"2afec80c",
   395 => x"fec80c58",
   396 => x"fec80c57",
   397 => x"fec80c84",
   398 => x"1a5a5376",
   399 => x"53848077",
   400 => x"25843884",
   401 => x"80537279",
   402 => x"24c4388c",
   403 => x"d904b5a8",
   404 => x"5185f32d",
   405 => x"72548cf5",
   406 => x"04bacc51",
   407 => x"99c82dfc",
   408 => x"80178119",
   409 => x"59578be4",
   410 => x"04820bfe",
   411 => x"c40c8154",
   412 => x"8cf50480",
   413 => x"5473baac",
   414 => x"0c02ac05",
   415 => x"0d0402f0",
   416 => x"050d7654",
   417 => x"a9b42d81",
   418 => x"f72d8151",
   419 => x"84e52d90",
   420 => x"53738338",
   421 => x"815372fe",
   422 => x"c40c840b",
   423 => x"fec40ca6",
   424 => x"ad2da6ad",
   425 => x"2d735275",
   426 => x"5189a02d",
   427 => x"b6e851ab",
   428 => x"922d8051",
   429 => x"84e52d02",
   430 => x"90050d04",
   431 => x"02f8050d",
   432 => x"80528251",
   433 => x"8cfe2d02",
   434 => x"88050d04",
   435 => x"02f8050d",
   436 => x"80528051",
   437 => x"8cfe2d02",
   438 => x"88050d04",
   439 => x"02f8050d",
   440 => x"81528051",
   441 => x"8cfe2d02",
   442 => x"88050d04",
   443 => x"02e8050d",
   444 => x"84b85187",
   445 => x"972d900b",
   446 => x"fec40c84",
   447 => x"b80bfec0",
   448 => x"0c840bfe",
   449 => x"c40c830b",
   450 => x"fecc0c81",
   451 => x"eef75188",
   452 => x"bf2d87f6",
   453 => x"2dbaac08",
   454 => x"fed40ca6",
   455 => x"c82da9a8",
   456 => x"2da6ad2d",
   457 => x"a6ad2d81",
   458 => x"f72d8151",
   459 => x"84e52da6",
   460 => x"ad2da6ad",
   461 => x"2d815184",
   462 => x"e52d8152",
   463 => x"815189a0",
   464 => x"2dbaac08",
   465 => x"802e8283",
   466 => x"38805184",
   467 => x"e52db6e8",
   468 => x"51ab922d",
   469 => x"bfb40853",
   470 => x"728b38bf",
   471 => x"b8085372",
   472 => x"802e818f",
   473 => x"38fed008",
   474 => x"70810651",
   475 => x"5372802e",
   476 => x"818138a9",
   477 => x"ae2dbfb4",
   478 => x"08bfb808",
   479 => x"555580ff",
   480 => x"75258438",
   481 => x"80ff5580",
   482 => x"ff742584",
   483 => x"3880ff54",
   484 => x"74ff8025",
   485 => x"8438ff80",
   486 => x"5573ff80",
   487 => x"258438ff",
   488 => x"8054bfb4",
   489 => x"08707631",
   490 => x"bfb40c53",
   491 => x"bfb80870",
   492 => x"7531bfb8",
   493 => x"0c53a9a8",
   494 => x"2db7a00b",
   495 => x"80f52d70",
   496 => x"812a7081",
   497 => x"06515456",
   498 => x"72802e89",
   499 => x"3874812c",
   500 => x"74812c55",
   501 => x"55758106",
   502 => x"5372802e",
   503 => x"85387381",
   504 => x"2c547488",
   505 => x"2b83fe80",
   506 => x"067481ff",
   507 => x"067107fe",
   508 => x"d00c53a7",
   509 => x"ad2daba2",
   510 => x"2dbaac08",
   511 => x"5486b52d",
   512 => x"baac08fe",
   513 => x"c00c87f6",
   514 => x"2dbaac08",
   515 => x"fed40c86",
   516 => x"b52dbaac",
   517 => x"08bac808",
   518 => x"2e9c38ba",
   519 => x"ac08bac8",
   520 => x"0c845373",
   521 => x"5184e52d",
   522 => x"a6ad2da6",
   523 => x"ad2dff13",
   524 => x"53728025",
   525 => x"ee387380",
   526 => x"2e89388a",
   527 => x"0bfec40c",
   528 => x"8ed40482",
   529 => x"0bfec40c",
   530 => x"8ed404b5",
   531 => x"b85185f3",
   532 => x"2d820bfe",
   533 => x"c40c800b",
   534 => x"baac0c02",
   535 => x"98050d04",
   536 => x"02e8050d",
   537 => x"77797b58",
   538 => x"55558053",
   539 => x"727625a3",
   540 => x"38747081",
   541 => x"055680f5",
   542 => x"2d747081",
   543 => x"055680f5",
   544 => x"2d525271",
   545 => x"712e8638",
   546 => x"81519195",
   547 => x"04811353",
   548 => x"90ec0480",
   549 => x"5170baac",
   550 => x"0c029805",
   551 => x"0d0402d8",
   552 => x"050d800b",
   553 => x"bee00cba",
   554 => x"d8528051",
   555 => x"a1bd2dba",
   556 => x"ac0854ba",
   557 => x"ac088c38",
   558 => x"b5d05185",
   559 => x"f32d7355",
   560 => x"96b90480",
   561 => x"56810bbf",
   562 => x"840c8853",
   563 => x"b5dc52bb",
   564 => x"8e5190e0",
   565 => x"2dbaac08",
   566 => x"762e0981",
   567 => x"068738ba",
   568 => x"ac08bf84",
   569 => x"0c8853b5",
   570 => x"e852bbaa",
   571 => x"5190e02d",
   572 => x"baac0887",
   573 => x"38baac08",
   574 => x"bf840cbf",
   575 => x"8408802e",
   576 => x"80f638be",
   577 => x"9e0b80f5",
   578 => x"2dbe9f0b",
   579 => x"80f52d71",
   580 => x"982b7190",
   581 => x"2b07bea0",
   582 => x"0b80f52d",
   583 => x"70882b72",
   584 => x"07bea10b",
   585 => x"80f52d71",
   586 => x"07bed60b",
   587 => x"80f52dbe",
   588 => x"d70b80f5",
   589 => x"2d71882b",
   590 => x"07535f54",
   591 => x"525a5657",
   592 => x"557381ab",
   593 => x"aa2e0981",
   594 => x"068d3875",
   595 => x"51a2df2d",
   596 => x"baac0856",
   597 => x"92e40473",
   598 => x"82d4d52e",
   599 => x"8738b5f4",
   600 => x"5193a504",
   601 => x"bad85275",
   602 => x"51a1bd2d",
   603 => x"baac0855",
   604 => x"baac0880",
   605 => x"2e83c238",
   606 => x"8853b5e8",
   607 => x"52bbaa51",
   608 => x"90e02dba",
   609 => x"ac088938",
   610 => x"810bbee0",
   611 => x"0c93ab04",
   612 => x"8853b5dc",
   613 => x"52bb8e51",
   614 => x"90e02dba",
   615 => x"ac08802e",
   616 => x"8a38b688",
   617 => x"5185f32d",
   618 => x"948504be",
   619 => x"d60b80f5",
   620 => x"2d547380",
   621 => x"d52e0981",
   622 => x"0680ca38",
   623 => x"bed70b80",
   624 => x"f52d5473",
   625 => x"81aa2e09",
   626 => x"8106ba38",
   627 => x"800bbad8",
   628 => x"0b80f52d",
   629 => x"56547481",
   630 => x"e92e8338",
   631 => x"81547481",
   632 => x"eb2e8c38",
   633 => x"80557375",
   634 => x"2e098106",
   635 => x"82cb38ba",
   636 => x"e30b80f5",
   637 => x"2d55748d",
   638 => x"38bae40b",
   639 => x"80f52d54",
   640 => x"73822e86",
   641 => x"38805596",
   642 => x"b904bae5",
   643 => x"0b80f52d",
   644 => x"70bed80c",
   645 => x"ff05bedc",
   646 => x"0cbae60b",
   647 => x"80f52dba",
   648 => x"e70b80f5",
   649 => x"2d587605",
   650 => x"77828029",
   651 => x"0570bee4",
   652 => x"0cbae80b",
   653 => x"80f52d70",
   654 => x"bef80cbe",
   655 => x"e0085957",
   656 => x"5876802e",
   657 => x"81a33888",
   658 => x"53b5e852",
   659 => x"bbaa5190",
   660 => x"e02dbaac",
   661 => x"0881e238",
   662 => x"bed80870",
   663 => x"842bbefc",
   664 => x"0c70bef4",
   665 => x"0cbafd0b",
   666 => x"80f52dba",
   667 => x"fc0b80f5",
   668 => x"2d718280",
   669 => x"2905bafe",
   670 => x"0b80f52d",
   671 => x"70848080",
   672 => x"2912baff",
   673 => x"0b80f52d",
   674 => x"7081800a",
   675 => x"291270bf",
   676 => x"800cbef8",
   677 => x"087129be",
   678 => x"e4080570",
   679 => x"bee80cbb",
   680 => x"850b80f5",
   681 => x"2dbb840b",
   682 => x"80f52d71",
   683 => x"82802905",
   684 => x"bb860b80",
   685 => x"f52d7084",
   686 => x"80802912",
   687 => x"bb870b80",
   688 => x"f52d7098",
   689 => x"2b81f00a",
   690 => x"06720570",
   691 => x"beec0cfe",
   692 => x"117e2977",
   693 => x"05bef00c",
   694 => x"52595243",
   695 => x"545e5152",
   696 => x"59525d57",
   697 => x"595796b7",
   698 => x"04baea0b",
   699 => x"80f52dba",
   700 => x"e90b80f5",
   701 => x"2d718280",
   702 => x"290570be",
   703 => x"fc0c70a0",
   704 => x"2983ff05",
   705 => x"70892a70",
   706 => x"bef40cba",
   707 => x"ef0b80f5",
   708 => x"2dbaee0b",
   709 => x"80f52d71",
   710 => x"82802905",
   711 => x"70bf800c",
   712 => x"7b71291e",
   713 => x"70bef00c",
   714 => x"7dbeec0c",
   715 => x"7305bee8",
   716 => x"0c555e51",
   717 => x"51555581",
   718 => x"5574baac",
   719 => x"0c02a805",
   720 => x"0d0402ec",
   721 => x"050d7670",
   722 => x"872c7180",
   723 => x"ff065556",
   724 => x"54bee008",
   725 => x"8a387388",
   726 => x"2c7481ff",
   727 => x"065455ba",
   728 => x"d852bee4",
   729 => x"081551a1",
   730 => x"bd2dbaac",
   731 => x"0854baac",
   732 => x"08802eb3",
   733 => x"38bee008",
   734 => x"802e9838",
   735 => x"728429ba",
   736 => x"d8057008",
   737 => x"5253a2df",
   738 => x"2dbaac08",
   739 => x"f00a0653",
   740 => x"97a50472",
   741 => x"10bad805",
   742 => x"7080e02d",
   743 => x"5253a38f",
   744 => x"2dbaac08",
   745 => x"53725473",
   746 => x"baac0c02",
   747 => x"94050d04",
   748 => x"02c8050d",
   749 => x"7f615f5b",
   750 => x"800bbeec",
   751 => x"08bef008",
   752 => x"595d56be",
   753 => x"e008762e",
   754 => x"8a38bed8",
   755 => x"08842b58",
   756 => x"97d904be",
   757 => x"f408842b",
   758 => x"58805978",
   759 => x"782781a9",
   760 => x"38788f06",
   761 => x"a0175754",
   762 => x"738f38ba",
   763 => x"d8527651",
   764 => x"811757a1",
   765 => x"bd2dbad8",
   766 => x"56807680",
   767 => x"f52d5654",
   768 => x"74742e83",
   769 => x"38815474",
   770 => x"81e52e80",
   771 => x"f6388170",
   772 => x"7506555d",
   773 => x"73802e80",
   774 => x"ea388b16",
   775 => x"80f52d98",
   776 => x"065a7980",
   777 => x"de388b53",
   778 => x"7d527551",
   779 => x"90e02dba",
   780 => x"ac0880cf",
   781 => x"389c1608",
   782 => x"51a2df2d",
   783 => x"baac0884",
   784 => x"1c0c9a16",
   785 => x"80e02d51",
   786 => x"a38f2dba",
   787 => x"ac08baac",
   788 => x"08881d0c",
   789 => x"baac0855",
   790 => x"55bee008",
   791 => x"802e9838",
   792 => x"941680e0",
   793 => x"2d51a38f",
   794 => x"2dbaac08",
   795 => x"902b83ff",
   796 => x"f00a0670",
   797 => x"16515473",
   798 => x"881c0c79",
   799 => x"7b0c7c54",
   800 => x"99bf0481",
   801 => x"195997db",
   802 => x"04bee008",
   803 => x"802eae38",
   804 => x"7b5196c2",
   805 => x"2dbaac08",
   806 => x"baac0880",
   807 => x"fffffff8",
   808 => x"06555c73",
   809 => x"80ffffff",
   810 => x"f82e9238",
   811 => x"baac08fe",
   812 => x"05bed808",
   813 => x"29bee808",
   814 => x"055797d9",
   815 => x"04805473",
   816 => x"baac0c02",
   817 => x"b8050d04",
   818 => x"02f4050d",
   819 => x"74700881",
   820 => x"05710c70",
   821 => x"08bedc08",
   822 => x"06535371",
   823 => x"8e388813",
   824 => x"085196c2",
   825 => x"2dbaac08",
   826 => x"88140c81",
   827 => x"0bbaac0c",
   828 => x"028c050d",
   829 => x"0402f005",
   830 => x"0d758811",
   831 => x"08fe05be",
   832 => x"d80829be",
   833 => x"e8081172",
   834 => x"08bedc08",
   835 => x"06057955",
   836 => x"535454a1",
   837 => x"bd2d0290",
   838 => x"050d0402",
   839 => x"f0050d75",
   840 => x"881108fe",
   841 => x"05bed808",
   842 => x"29bee808",
   843 => x"117208be",
   844 => x"dc080605",
   845 => x"79555354",
   846 => x"549ffd2d",
   847 => x"0290050d",
   848 => x"04bee008",
   849 => x"baac0c04",
   850 => x"02f4050d",
   851 => x"d45281ff",
   852 => x"720c7108",
   853 => x"5381ff72",
   854 => x"0c72882b",
   855 => x"83fe8006",
   856 => x"72087081",
   857 => x"ff065152",
   858 => x"5381ff72",
   859 => x"0c727107",
   860 => x"882b7208",
   861 => x"7081ff06",
   862 => x"51525381",
   863 => x"ff720c72",
   864 => x"7107882b",
   865 => x"72087081",
   866 => x"ff067207",
   867 => x"baac0c52",
   868 => x"53028c05",
   869 => x"0d0402f4",
   870 => x"050d7476",
   871 => x"7181ff06",
   872 => x"d40c5353",
   873 => x"bf880885",
   874 => x"3871892b",
   875 => x"5271982a",
   876 => x"d40c7190",
   877 => x"2a7081ff",
   878 => x"06d40c51",
   879 => x"71882a70",
   880 => x"81ff06d4",
   881 => x"0c517181",
   882 => x"ff06d40c",
   883 => x"72902a70",
   884 => x"81ff06d4",
   885 => x"0c51d408",
   886 => x"7081ff06",
   887 => x"515182b8",
   888 => x"bf527081",
   889 => x"ff2e0981",
   890 => x"06943881",
   891 => x"ff0bd40c",
   892 => x"d4087081",
   893 => x"ff06ff14",
   894 => x"54515171",
   895 => x"e53870ba",
   896 => x"ac0c028c",
   897 => x"050d0402",
   898 => x"fc050d81",
   899 => x"c75181ff",
   900 => x"0bd40cff",
   901 => x"11517080",
   902 => x"25f43802",
   903 => x"84050d04",
   904 => x"02f0050d",
   905 => x"9c872d8f",
   906 => x"cf538052",
   907 => x"87fc80f7",
   908 => x"519b962d",
   909 => x"baac0854",
   910 => x"baac0881",
   911 => x"2e098106",
   912 => x"a33881ff",
   913 => x"0bd40c82",
   914 => x"0a52849c",
   915 => x"80e9519b",
   916 => x"962dbaac",
   917 => x"088b3881",
   918 => x"ff0bd40c",
   919 => x"73539cea",
   920 => x"049c872d",
   921 => x"ff135372",
   922 => x"c13872ba",
   923 => x"ac0c0290",
   924 => x"050d0402",
   925 => x"f4050d81",
   926 => x"ff0bd40c",
   927 => x"93538052",
   928 => x"87fc80c1",
   929 => x"519b962d",
   930 => x"baac088b",
   931 => x"3881ff0b",
   932 => x"d40c8153",
   933 => x"9da0049c",
   934 => x"872dff13",
   935 => x"5372df38",
   936 => x"72baac0c",
   937 => x"028c050d",
   938 => x"0402f005",
   939 => x"0d9c872d",
   940 => x"83aa5284",
   941 => x"9c80c851",
   942 => x"9b962dba",
   943 => x"ac08812e",
   944 => x"09810692",
   945 => x"389ac82d",
   946 => x"baac0883",
   947 => x"ffff0653",
   948 => x"7283aa2e",
   949 => x"97389cf3",
   950 => x"2d9de704",
   951 => x"81549ecc",
   952 => x"04b69451",
   953 => x"85f32d80",
   954 => x"549ecc04",
   955 => x"81ff0bd4",
   956 => x"0cb1539c",
   957 => x"a02dbaac",
   958 => x"08802e80",
   959 => x"c0388052",
   960 => x"87fc80fa",
   961 => x"519b962d",
   962 => x"baac08b1",
   963 => x"3881ff0b",
   964 => x"d40cd408",
   965 => x"5381ff0b",
   966 => x"d40c81ff",
   967 => x"0bd40c81",
   968 => x"ff0bd40c",
   969 => x"81ff0bd4",
   970 => x"0c72862a",
   971 => x"708106ba",
   972 => x"ac085651",
   973 => x"5372802e",
   974 => x"93389ddc",
   975 => x"0472822e",
   976 => x"ff9f38ff",
   977 => x"135372ff",
   978 => x"aa387254",
   979 => x"73baac0c",
   980 => x"0290050d",
   981 => x"0402f005",
   982 => x"0d810bbf",
   983 => x"880c8454",
   984 => x"d008708f",
   985 => x"2a708106",
   986 => x"51515372",
   987 => x"f33872d0",
   988 => x"0c9c872d",
   989 => x"b6a45185",
   990 => x"f32dd008",
   991 => x"708f2a70",
   992 => x"81065151",
   993 => x"5372f338",
   994 => x"810bd00c",
   995 => x"b1538052",
   996 => x"84d480c0",
   997 => x"519b962d",
   998 => x"baac0881",
   999 => x"2ea13872",
  1000 => x"822e0981",
  1001 => x"068c38b6",
  1002 => x"b05185f3",
  1003 => x"2d80539f",
  1004 => x"f404ff13",
  1005 => x"5372d738",
  1006 => x"ff145473",
  1007 => x"ffa2389d",
  1008 => x"a92dbaac",
  1009 => x"08bf880c",
  1010 => x"baac088b",
  1011 => x"38815287",
  1012 => x"fc80d051",
  1013 => x"9b962d81",
  1014 => x"ff0bd40c",
  1015 => x"d008708f",
  1016 => x"2a708106",
  1017 => x"51515372",
  1018 => x"f33872d0",
  1019 => x"0c81ff0b",
  1020 => x"d40c8153",
  1021 => x"72baac0c",
  1022 => x"0290050d",
  1023 => x"0402e805",
  1024 => x"0d785681",
  1025 => x"ff0bd40c",
  1026 => x"d008708f",
  1027 => x"2a708106",
  1028 => x"51515372",
  1029 => x"f3388281",
  1030 => x"0bd00c81",
  1031 => x"ff0bd40c",
  1032 => x"775287fc",
  1033 => x"80d8519b",
  1034 => x"962dbaac",
  1035 => x"08802e8c",
  1036 => x"38b6c851",
  1037 => x"85f32d81",
  1038 => x"53a1b404",
  1039 => x"81ff0bd4",
  1040 => x"0c81fe0b",
  1041 => x"d40c80ff",
  1042 => x"55757084",
  1043 => x"05570870",
  1044 => x"982ad40c",
  1045 => x"70902c70",
  1046 => x"81ff06d4",
  1047 => x"0c547088",
  1048 => x"2c7081ff",
  1049 => x"06d40c54",
  1050 => x"7081ff06",
  1051 => x"d40c54ff",
  1052 => x"15557480",
  1053 => x"25d33881",
  1054 => x"ff0bd40c",
  1055 => x"81ff0bd4",
  1056 => x"0c81ff0b",
  1057 => x"d40c868d",
  1058 => x"a05481ff",
  1059 => x"0bd40cd4",
  1060 => x"0881ff06",
  1061 => x"55748738",
  1062 => x"ff145473",
  1063 => x"ed3881ff",
  1064 => x"0bd40cd0",
  1065 => x"08708f2a",
  1066 => x"70810651",
  1067 => x"515372f3",
  1068 => x"3872d00c",
  1069 => x"72baac0c",
  1070 => x"0298050d",
  1071 => x"0402e805",
  1072 => x"0d785580",
  1073 => x"5681ff0b",
  1074 => x"d40cd008",
  1075 => x"708f2a70",
  1076 => x"81065151",
  1077 => x"5372f338",
  1078 => x"82810bd0",
  1079 => x"0c81ff0b",
  1080 => x"d40c7752",
  1081 => x"87fc80d1",
  1082 => x"519b962d",
  1083 => x"80dbc6df",
  1084 => x"54baac08",
  1085 => x"802e8a38",
  1086 => x"b5a85185",
  1087 => x"f32da2cf",
  1088 => x"0481ff0b",
  1089 => x"d40cd408",
  1090 => x"7081ff06",
  1091 => x"51537281",
  1092 => x"fe2e0981",
  1093 => x"069d3880",
  1094 => x"ff539ac8",
  1095 => x"2dbaac08",
  1096 => x"75708405",
  1097 => x"570cff13",
  1098 => x"53728025",
  1099 => x"ed388156",
  1100 => x"a2b904ff",
  1101 => x"145473c9",
  1102 => x"3881ff0b",
  1103 => x"d40cd008",
  1104 => x"708f2a70",
  1105 => x"81065151",
  1106 => x"5372f338",
  1107 => x"72d00c75",
  1108 => x"baac0c02",
  1109 => x"98050d04",
  1110 => x"bf8808ba",
  1111 => x"ac0c0402",
  1112 => x"f4050d74",
  1113 => x"70882a83",
  1114 => x"fe800670",
  1115 => x"72982a07",
  1116 => x"72882b87",
  1117 => x"fc808006",
  1118 => x"73982b81",
  1119 => x"f00a0671",
  1120 => x"730707ba",
  1121 => x"ac0c5651",
  1122 => x"5351028c",
  1123 => x"050d0402",
  1124 => x"f8050d02",
  1125 => x"8e0580f5",
  1126 => x"2d74882b",
  1127 => x"077083ff",
  1128 => x"ff06baac",
  1129 => x"0c510288",
  1130 => x"050d0402",
  1131 => x"fc050d72",
  1132 => x"5180710c",
  1133 => x"800b8412",
  1134 => x"0c028405",
  1135 => x"0d0402f0",
  1136 => x"050d7570",
  1137 => x"08841208",
  1138 => x"535353ff",
  1139 => x"5471712e",
  1140 => x"a838a9ae",
  1141 => x"2d841308",
  1142 => x"70842914",
  1143 => x"88117008",
  1144 => x"7081ff06",
  1145 => x"84180881",
  1146 => x"11870684",
  1147 => x"1a0c5351",
  1148 => x"55515151",
  1149 => x"a9a82d71",
  1150 => x"5473baac",
  1151 => x"0c029005",
  1152 => x"0d0402f4",
  1153 => x"050da9ae",
  1154 => x"2de008e4",
  1155 => x"08718b2a",
  1156 => x"70810651",
  1157 => x"53545270",
  1158 => x"802e9d38",
  1159 => x"bf8c0870",
  1160 => x"8429bf94",
  1161 => x"057381ff",
  1162 => x"06710c51",
  1163 => x"51bf8c08",
  1164 => x"81118706",
  1165 => x"bf8c0c51",
  1166 => x"728b2a70",
  1167 => x"81065151",
  1168 => x"70802e81",
  1169 => x"9b38b9dc",
  1170 => x"088429bf",
  1171 => x"c0057381",
  1172 => x"ff06710c",
  1173 => x"51b9dc08",
  1174 => x"8105b9dc",
  1175 => x"0c850bb9",
  1176 => x"d80cb9dc",
  1177 => x"08b9d408",
  1178 => x"2e098106",
  1179 => x"81af3880",
  1180 => x"0bb9dc0c",
  1181 => x"bfd00881",
  1182 => x"a438bfc0",
  1183 => x"08700970",
  1184 => x"8306fecc",
  1185 => x"0c527085",
  1186 => x"2a708106",
  1187 => x"51525270",
  1188 => x"802e9038",
  1189 => x"bfb808bf",
  1190 => x"c808fe80",
  1191 => x"32115151",
  1192 => x"a5ac04bf",
  1193 => x"b808bfc8",
  1194 => x"08115151",
  1195 => x"70bfb80c",
  1196 => x"71842a70",
  1197 => x"81065151",
  1198 => x"70802e93",
  1199 => x"38bfb408",
  1200 => x"bfc40881",
  1201 => x"ff321181",
  1202 => x"11515151",
  1203 => x"a5d904bf",
  1204 => x"b40870bf",
  1205 => x"c4083151",
  1206 => x"5170bfb4",
  1207 => x"0ca69d04",
  1208 => x"b9d808ff",
  1209 => x"05b9d80c",
  1210 => x"b9d808ff",
  1211 => x"2e098106",
  1212 => x"ac38b9dc",
  1213 => x"08802e92",
  1214 => x"38810bbf",
  1215 => x"d00c870b",
  1216 => x"b9d40831",
  1217 => x"b9d40ca6",
  1218 => x"9804bfd0",
  1219 => x"08517080",
  1220 => x"2e8638ff",
  1221 => x"11bfd00c",
  1222 => x"800bb9dc",
  1223 => x"0c800bbf",
  1224 => x"bc0ca9a1",
  1225 => x"2da9a82d",
  1226 => x"028c050d",
  1227 => x"0402fc05",
  1228 => x"0da9ae2d",
  1229 => x"810bbfbc",
  1230 => x"0ca9a82d",
  1231 => x"bfbc0851",
  1232 => x"70fa3802",
  1233 => x"84050d04",
  1234 => x"02f8050d",
  1235 => x"bf8c51a3",
  1236 => x"ab2d800b",
  1237 => x"bfd00c83",
  1238 => x"0bb9d40c",
  1239 => x"e408708c",
  1240 => x"2a708106",
  1241 => x"51515271",
  1242 => x"802e8638",
  1243 => x"840bb9d4",
  1244 => x"0ce40870",
  1245 => x"8d2a7081",
  1246 => x"06515152",
  1247 => x"71802e9f",
  1248 => x"38870bb9",
  1249 => x"d40831b9",
  1250 => x"d40ce408",
  1251 => x"708a2a70",
  1252 => x"81065151",
  1253 => x"5271802e",
  1254 => x"f13881f4",
  1255 => x"0be40ca4",
  1256 => x"8251a99d",
  1257 => x"2da8c72d",
  1258 => x"0288050d",
  1259 => x"0402f405",
  1260 => x"0da8af04",
  1261 => x"baac0881",
  1262 => x"f02e0981",
  1263 => x"06893881",
  1264 => x"0bbaa00c",
  1265 => x"a8af04ba",
  1266 => x"ac0881e0",
  1267 => x"2e098106",
  1268 => x"8938810b",
  1269 => x"baa40ca8",
  1270 => x"af04baac",
  1271 => x"0852baa4",
  1272 => x"08802e88",
  1273 => x"38baac08",
  1274 => x"81800552",
  1275 => x"71842c72",
  1276 => x"8f065353",
  1277 => x"baa00880",
  1278 => x"2e993872",
  1279 => x"8429b9e0",
  1280 => x"05721381",
  1281 => x"712b7009",
  1282 => x"73080673",
  1283 => x"0c515353",
  1284 => x"a8a50472",
  1285 => x"8429b9e0",
  1286 => x"05721383",
  1287 => x"712b7208",
  1288 => x"07720c53",
  1289 => x"53800bba",
  1290 => x"a40c800b",
  1291 => x"baa00cbf",
  1292 => x"8c51a3be",
  1293 => x"2dbaac08",
  1294 => x"ff24fef8",
  1295 => x"38800bba",
  1296 => x"ac0c028c",
  1297 => x"050d0402",
  1298 => x"f8050db9",
  1299 => x"e0528f51",
  1300 => x"80727084",
  1301 => x"05540cff",
  1302 => x"11517080",
  1303 => x"25f23802",
  1304 => x"88050d04",
  1305 => x"02f0050d",
  1306 => x"7551a9ae",
  1307 => x"2d70822c",
  1308 => x"fc06b9e0",
  1309 => x"1172109e",
  1310 => x"06710870",
  1311 => x"722a7083",
  1312 => x"0682742b",
  1313 => x"70097406",
  1314 => x"760c5451",
  1315 => x"56575351",
  1316 => x"53a9a82d",
  1317 => x"71baac0c",
  1318 => x"0290050d",
  1319 => x"0471980c",
  1320 => x"04ffb008",
  1321 => x"baac0c04",
  1322 => x"810bffb0",
  1323 => x"0c04800b",
  1324 => x"ffb00c04",
  1325 => x"02fc050d",
  1326 => x"800bbaa8",
  1327 => x"0c805184",
  1328 => x"e52d0284",
  1329 => x"050d0402",
  1330 => x"ec050d76",
  1331 => x"54805287",
  1332 => x"0b881580",
  1333 => x"f52d5653",
  1334 => x"74722483",
  1335 => x"38a05372",
  1336 => x"5182ee2d",
  1337 => x"81128b15",
  1338 => x"80f52d54",
  1339 => x"52727225",
  1340 => x"de380294",
  1341 => x"050d0402",
  1342 => x"f0050dbf",
  1343 => x"d8085481",
  1344 => x"f72d800b",
  1345 => x"bfdc0c73",
  1346 => x"08802e81",
  1347 => x"8038820b",
  1348 => x"bac00cbf",
  1349 => x"dc088f06",
  1350 => x"babc0c73",
  1351 => x"08527183",
  1352 => x"2e963871",
  1353 => x"83268938",
  1354 => x"71812eaf",
  1355 => x"38aaf804",
  1356 => x"71852e9f",
  1357 => x"38aaf804",
  1358 => x"881480f5",
  1359 => x"2d841508",
  1360 => x"b6d85354",
  1361 => x"5285f32d",
  1362 => x"71842913",
  1363 => x"70085252",
  1364 => x"aafc0473",
  1365 => x"51a9c72d",
  1366 => x"aaf804bf",
  1367 => x"d4088815",
  1368 => x"082c7081",
  1369 => x"06515271",
  1370 => x"802e8738",
  1371 => x"b6dc51aa",
  1372 => x"f504b6e0",
  1373 => x"5185f32d",
  1374 => x"84140851",
  1375 => x"85f32dbf",
  1376 => x"dc088105",
  1377 => x"bfdc0c8c",
  1378 => x"1454aa87",
  1379 => x"04029005",
  1380 => x"0d0471bf",
  1381 => x"d80ca9f7",
  1382 => x"2dbfdc08",
  1383 => x"ff05bfe0",
  1384 => x"0c0402e8",
  1385 => x"050d800b",
  1386 => x"bfd80856",
  1387 => x"5680f851",
  1388 => x"a8e42dba",
  1389 => x"ac08812a",
  1390 => x"70810651",
  1391 => x"5271762e",
  1392 => x"0981069b",
  1393 => x"388751a8",
  1394 => x"e42dbaac",
  1395 => x"08812a70",
  1396 => x"81065152",
  1397 => x"71762eba",
  1398 => x"38abdf04",
  1399 => x"a7ad2d87",
  1400 => x"51a8e42d",
  1401 => x"baac08f4",
  1402 => x"38abef04",
  1403 => x"a7ad2d80",
  1404 => x"f851a8e4",
  1405 => x"2dbaac08",
  1406 => x"f338baa8",
  1407 => x"08813270",
  1408 => x"baa80c70",
  1409 => x"525284e5",
  1410 => x"2dbaa808",
  1411 => x"802e8338",
  1412 => x"8156baa8",
  1413 => x"08a23880",
  1414 => x"da51a8e4",
  1415 => x"2d81f551",
  1416 => x"a8e42d81",
  1417 => x"f251a8e4",
  1418 => x"2d81eb51",
  1419 => x"a8e42d81",
  1420 => x"f451a8e4",
  1421 => x"2db08c04",
  1422 => x"81f551a8",
  1423 => x"e42dbaac",
  1424 => x"08812a70",
  1425 => x"81065152",
  1426 => x"71802e91",
  1427 => x"38bfe008",
  1428 => x"5271802e",
  1429 => x"8838ff12",
  1430 => x"bfe00c81",
  1431 => x"5681f251",
  1432 => x"a8e42dba",
  1433 => x"ac08812a",
  1434 => x"70810651",
  1435 => x"5271802e",
  1436 => x"9738bfdc",
  1437 => x"08ff05bf",
  1438 => x"e0085452",
  1439 => x"72722588",
  1440 => x"388113bf",
  1441 => x"e00c8156",
  1442 => x"bfe00870",
  1443 => x"53547380",
  1444 => x"2e8a388c",
  1445 => x"15ff1555",
  1446 => x"55ad8e04",
  1447 => x"820bbac0",
  1448 => x"0c718f06",
  1449 => x"babc0c81",
  1450 => x"eb51a8e4",
  1451 => x"2dbaac08",
  1452 => x"812a7081",
  1453 => x"06515271",
  1454 => x"802eaf38",
  1455 => x"81567408",
  1456 => x"852e0981",
  1457 => x"06a43888",
  1458 => x"1580f52d",
  1459 => x"ff055271",
  1460 => x"881681b7",
  1461 => x"2d71982b",
  1462 => x"52718025",
  1463 => x"8838800b",
  1464 => x"881681b7",
  1465 => x"2d7451a9",
  1466 => x"c72d81f4",
  1467 => x"51a8e42d",
  1468 => x"baac0881",
  1469 => x"2a708106",
  1470 => x"51527180",
  1471 => x"2eb53881",
  1472 => x"56740885",
  1473 => x"2e098106",
  1474 => x"aa388815",
  1475 => x"80f52d76",
  1476 => x"05527188",
  1477 => x"1681b72d",
  1478 => x"7181ff06",
  1479 => x"8b1680f5",
  1480 => x"2d545272",
  1481 => x"72278738",
  1482 => x"72881681",
  1483 => x"b72d7451",
  1484 => x"a9c72d80",
  1485 => x"da51a8e4",
  1486 => x"2dbaac08",
  1487 => x"812a7081",
  1488 => x"06515271",
  1489 => x"802e80fe",
  1490 => x"38bfd808",
  1491 => x"bfe00855",
  1492 => x"5373802e",
  1493 => x"8a388c13",
  1494 => x"ff155553",
  1495 => x"aed10472",
  1496 => x"08527182",
  1497 => x"2ea63871",
  1498 => x"82268938",
  1499 => x"71812ea5",
  1500 => x"38afcb04",
  1501 => x"71832ead",
  1502 => x"3871842e",
  1503 => x"09810680",
  1504 => x"ca388813",
  1505 => x"0851ab92",
  1506 => x"2dafcb04",
  1507 => x"88130852",
  1508 => x"712dafcb",
  1509 => x"04810b88",
  1510 => x"14082bbf",
  1511 => x"d40832bf",
  1512 => x"d40cafc0",
  1513 => x"04881380",
  1514 => x"f52d8105",
  1515 => x"8b1480f5",
  1516 => x"2d535471",
  1517 => x"74248338",
  1518 => x"80547388",
  1519 => x"1481b72d",
  1520 => x"a9f72daf",
  1521 => x"cb047580",
  1522 => x"2ebe3880",
  1523 => x"54800bba",
  1524 => x"c00c738f",
  1525 => x"06babc0c",
  1526 => x"a05273bf",
  1527 => x"e0082e09",
  1528 => x"81069838",
  1529 => x"bfdc08ff",
  1530 => x"05743270",
  1531 => x"09810570",
  1532 => x"72079f2a",
  1533 => x"91713151",
  1534 => x"51535371",
  1535 => x"5182ee2d",
  1536 => x"8114548e",
  1537 => x"7425c638",
  1538 => x"baa80852",
  1539 => x"71baac0c",
  1540 => x"0298050d",
  1541 => x"04000000",
  1542 => x"00ffffff",
  1543 => x"ff00ffff",
  1544 => x"ffff00ff",
  1545 => x"ffffff00",
  1546 => x"4f707469",
  1547 => x"6f6e7320",
  1548 => x"10000000",
  1549 => x"536f756e",
  1550 => x"64201000",
  1551 => x"54757262",
  1552 => x"6f000000",
  1553 => x"4d6f7573",
  1554 => x"6520456d",
  1555 => x"756c6174",
  1556 => x"696f6e00",
  1557 => x"53617665",
  1558 => x"20616e64",
  1559 => x"20526573",
  1560 => x"65740000",
  1561 => x"48617264",
  1562 => x"20526573",
  1563 => x"65740000",
  1564 => x"52657365",
  1565 => x"74000000",
  1566 => x"45786974",
  1567 => x"00000000",
  1568 => x"20205363",
  1569 => x"616c696e",
  1570 => x"6720313a",
  1571 => x"31000000",
  1572 => x"20205363",
  1573 => x"616c696e",
  1574 => x"6720323a",
  1575 => x"31000000",
  1576 => x"20205363",
  1577 => x"616c696e",
  1578 => x"6720323a",
  1579 => x"32000000",
  1580 => x"20205363",
  1581 => x"616c696e",
  1582 => x"6720343a",
  1583 => x"32000000",
  1584 => x"4d617374",
  1585 => x"65720000",
  1586 => x"4f504c4c",
  1587 => x"00000000",
  1588 => x"53434300",
  1589 => x"50534700",
  1590 => x"4261636b",
  1591 => x"00000000",
  1592 => x"5363616e",
  1593 => x"6c696e65",
  1594 => x"73000000",
  1595 => x"53442043",
  1596 => x"61726400",
  1597 => x"4a617061",
  1598 => x"6e657365",
  1599 => x"206b6579",
  1600 => x"206c6179",
  1601 => x"6f757400",
  1602 => x"32303438",
  1603 => x"4b422052",
  1604 => x"414d0000",
  1605 => x"34303936",
  1606 => x"4b422052",
  1607 => x"414d0000",
  1608 => x"536c323a",
  1609 => x"204e6f6e",
  1610 => x"65000000",
  1611 => x"536c323a",
  1612 => x"20455345",
  1613 => x"2d52414d",
  1614 => x"20314d42",
  1615 => x"2f415343",
  1616 => x"49493800",
  1617 => x"536c323a",
  1618 => x"20455345",
  1619 => x"2d534343",
  1620 => x"20314d42",
  1621 => x"2f534343",
  1622 => x"2d490000",
  1623 => x"536c323a",
  1624 => x"20455345",
  1625 => x"2d52414d",
  1626 => x"20314d42",
  1627 => x"2f415343",
  1628 => x"49493136",
  1629 => x"00000000",
  1630 => x"536c313a",
  1631 => x"204e6f6e",
  1632 => x"65000000",
  1633 => x"536c313a",
  1634 => x"20455345",
  1635 => x"2d534343",
  1636 => x"20314d42",
  1637 => x"2f534343",
  1638 => x"2d490000",
  1639 => x"536c313a",
  1640 => x"204d6567",
  1641 => x"6152414d",
  1642 => x"00000000",
  1643 => x"56474120",
  1644 => x"2d203331",
  1645 => x"4b487a2c",
  1646 => x"20363048",
  1647 => x"7a000000",
  1648 => x"56474120",
  1649 => x"2d203331",
  1650 => x"4b487a2c",
  1651 => x"20353048",
  1652 => x"7a000000",
  1653 => x"5456202d",
  1654 => x"20343830",
  1655 => x"692c2036",
  1656 => x"30487a00",
  1657 => x"496e6974",
  1658 => x"69616c69",
  1659 => x"7a696e67",
  1660 => x"20534420",
  1661 => x"63617264",
  1662 => x"0a000000",
  1663 => x"53444843",
  1664 => x"206e6f74",
  1665 => x"20737570",
  1666 => x"706f7274",
  1667 => x"65643b00",
  1668 => x"46617433",
  1669 => x"32206e6f",
  1670 => x"74207375",
  1671 => x"70706f72",
  1672 => x"7465643b",
  1673 => x"00000000",
  1674 => x"0a646973",
  1675 => x"61626c69",
  1676 => x"6e672053",
  1677 => x"44206361",
  1678 => x"72640a10",
  1679 => x"204f4b0a",
  1680 => x"00000000",
  1681 => x"4f434d53",
  1682 => x"58202020",
  1683 => x"43464700",
  1684 => x"54727969",
  1685 => x"6e67204d",
  1686 => x"53583342",
  1687 => x"494f532e",
  1688 => x"5359530a",
  1689 => x"00000000",
  1690 => x"4d535833",
  1691 => x"42494f53",
  1692 => x"53595300",
  1693 => x"54727969",
  1694 => x"6e672042",
  1695 => x"494f535f",
  1696 => x"4d32502e",
  1697 => x"524f4d0a",
  1698 => x"00000000",
  1699 => x"42494f53",
  1700 => x"5f4d3250",
  1701 => x"524f4d00",
  1702 => x"4c6f6164",
  1703 => x"696e6720",
  1704 => x"42494f53",
  1705 => x"0a000000",
  1706 => x"52656164",
  1707 => x"20666169",
  1708 => x"6c65640a",
  1709 => x"00000000",
  1710 => x"4c6f6164",
  1711 => x"696e6720",
  1712 => x"42494f53",
  1713 => x"20666169",
  1714 => x"6c65640a",
  1715 => x"00000000",
  1716 => x"4d425220",
  1717 => x"6661696c",
  1718 => x"0a000000",
  1719 => x"46415431",
  1720 => x"36202020",
  1721 => x"00000000",
  1722 => x"46415433",
  1723 => x"32202020",
  1724 => x"00000000",
  1725 => x"4e6f2070",
  1726 => x"61727469",
  1727 => x"74696f6e",
  1728 => x"20736967",
  1729 => x"0a000000",
  1730 => x"42616420",
  1731 => x"70617274",
  1732 => x"0a000000",
  1733 => x"53444843",
  1734 => x"20657272",
  1735 => x"6f72210a",
  1736 => x"00000000",
  1737 => x"53442069",
  1738 => x"6e69742e",
  1739 => x"2e2e0a00",
  1740 => x"53442063",
  1741 => x"61726420",
  1742 => x"72657365",
  1743 => x"74206661",
  1744 => x"696c6564",
  1745 => x"210a0000",
  1746 => x"57726974",
  1747 => x"65206661",
  1748 => x"696c6564",
  1749 => x"0a000000",
  1750 => x"16200000",
  1751 => x"14200000",
  1752 => x"15200000",
  1753 => x"00000002",
  1754 => x"00000004",
  1755 => x"00001828",
  1756 => x"00001c38",
  1757 => x"00000004",
  1758 => x"00001834",
  1759 => x"00001bf0",
  1760 => x"00000001",
  1761 => x"0000183c",
  1762 => x"00000007",
  1763 => x"00000001",
  1764 => x"00001844",
  1765 => x"0000000a",
  1766 => x"00000003",
  1767 => x"00001be0",
  1768 => x"00000004",
  1769 => x"00000002",
  1770 => x"00001854",
  1771 => x"000006bc",
  1772 => x"00000002",
  1773 => x"00001864",
  1774 => x"000006dc",
  1775 => x"00000002",
  1776 => x"00001870",
  1777 => x"000006cc",
  1778 => x"00000002",
  1779 => x"00001878",
  1780 => x"000014b4",
  1781 => x"00000000",
  1782 => x"00000000",
  1783 => x"00000000",
  1784 => x"00001880",
  1785 => x"00001890",
  1786 => x"000018a0",
  1787 => x"000018b0",
  1788 => x"00000005",
  1789 => x"000018c0",
  1790 => x"00000007",
  1791 => x"00000005",
  1792 => x"000018c8",
  1793 => x"00000007",
  1794 => x"00000005",
  1795 => x"000018d0",
  1796 => x"00000007",
  1797 => x"00000005",
  1798 => x"000018d4",
  1799 => x"00000007",
  1800 => x"00000004",
  1801 => x"000018d8",
  1802 => x"00001b68",
  1803 => x"00000000",
  1804 => x"00000000",
  1805 => x"00000000",
  1806 => x"00000003",
  1807 => x"00001cc8",
  1808 => x"00000003",
  1809 => x"00000001",
  1810 => x"000018e0",
  1811 => x"0000000b",
  1812 => x"00000001",
  1813 => x"000018ec",
  1814 => x"00000002",
  1815 => x"00000003",
  1816 => x"00001cbc",
  1817 => x"00000003",
  1818 => x"00000003",
  1819 => x"00001cac",
  1820 => x"00000004",
  1821 => x"00000001",
  1822 => x"000018f4",
  1823 => x"00000006",
  1824 => x"00000003",
  1825 => x"00001ca4",
  1826 => x"00000002",
  1827 => x"00000004",
  1828 => x"000018d8",
  1829 => x"00001b68",
  1830 => x"00000000",
  1831 => x"00000000",
  1832 => x"00000000",
  1833 => x"00001908",
  1834 => x"00001914",
  1835 => x"00001920",
  1836 => x"0000192c",
  1837 => x"00001944",
  1838 => x"0000195c",
  1839 => x"00001978",
  1840 => x"00001984",
  1841 => x"0000199c",
  1842 => x"000019ac",
  1843 => x"000019c0",
  1844 => x"000019d4",
  1845 => x"00000003",
  1846 => x"00000000",
  1847 => x"00000000",
  1848 => x"00000000",
  1849 => x"00000000",
  1850 => x"00000000",
  1851 => x"00000000",
  1852 => x"00000000",
  1853 => x"00000000",
  1854 => x"00000000",
  1855 => x"00000000",
  1856 => x"00000000",
  1857 => x"00000000",
  1858 => x"00000000",
  1859 => x"00000000",
  1860 => x"00000000",
  1861 => x"00000000",
  1862 => x"00000000",
  1863 => x"00000000",
  1864 => x"00000000",
  1865 => x"00000000",
  1866 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

